* NGSPICE file created from raven.ext - technology: EFXH018D

* Need include to schematic netlist for CORNERESDF
* Unknown black-box entry CORNERESDF
.subckt CORNERESDF GNDR VDDR VDD VDDO GNDO

* Need include to schematic netlist for FILLER01F
* Unknown black-box entry FILLER01F
.subckt FILLER01F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for FILLER10F
* Unknown black-box entry FILLER10F
.subckt FILLER10F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for FILLER20F
* Unknown black-box entry FILLER20F
.subckt FILLER20F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for FILLER50F
* Unknown black-box entry FILLER50F
.subckt FILLER50F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for VDDPADF
* Unknown black-box entry VDDPADF
.subckt VDDPADF VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for VDDORPADF
* Unknown black-box entry VDDORPADF
.subckt VDDORPADF VDDOR GNDR GNDO VDD

* Need include to schematic netlist for GNDORPADF
* Unknown black-box entry GNDORPADF
.subckt GNDORPADF VDDO VDDR VDD GNDOR

* Need include to schematic netlist for ICF
* Unknown black-box entry ICF
.subckt ICF PO PI Y PAD VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for BT4F
* Unknown black-box entry BT4F
.subckt BT4F EN A PAD VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for BBC4F
* Unknown black-box entry BBC4F
.subckt BBC4F EN A Y PO PI PAD VDDO GNDO GNDR VDDR VDD

* Need include to schematic netlist for FILLER40F
* Unknown black-box entry FILLER40F
.subckt FILLER40F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for POWERCUTVDD3FC
* Unknown black-box entry POWERCUTVDD3FC
.subckt POWERCUTVDD3FC VDDO VDDR GNDR GNDO

* Need include to schematic netlist for VDDPADFC
* Unknown black-box entry VDDPADFC
.subckt VDDPADFC VDDO VDDR GNDR GNDO VDD3

* Need include to schematic netlist for BT4FC
* Unknown black-box entry BT4FC
.subckt BT4FC EN A PAD VDDO VDDR GNDR GNDO VDD3

* Need include to schematic netlist for ICFC
* Unknown black-box entry ICFC
.subckt ICFC PO PI Y PAD VDDO VDDR GNDR GNDO VDD3

* Need include to schematic netlist for FILLER20FC
* Unknown black-box entry FILLER20FC
.subckt FILLER20FC VDDO VDDR GNDR GNDO VDD3

* Need include to schematic netlist for BBCUD4F
* Unknown black-box entry BBCUD4F
.subckt BBCUD4F EN A Y PO PI PUEN PDEN PAD VDDO GNDO GNDR VDDR VDD

* Need include to schematic netlist for APR00DF
* Unknown black-box entry APR00DF
.subckt APR00DF PAD VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for aregc01_3v3
* Unknown black-box entry aregc01_3v3
.subckt aregc01_3v3 OUT EN VIN3 ENB VDD VDDR GNDR GNDO VDDO

* Need include to schematic netlist for FILLER02F
* Unknown black-box entry FILLER02F
.subckt FILLER02F VDDO VDDR GNDR GNDO VDD

* Need include to schematic netlist for axtoc02_3v3
* Unknown black-box entry axtoc02_3v3
.subckt axtoc02_3v3 GNDO VDDO GNDR VDDR VDD XI XO CLK EN

.subckt raven_padframe VDD3V3 VDD1V8 BBCUD4F_0|PI BBCUD4F_4|EN gpio<10> VDD1V8 VDD3V3  XCLK comp_inn BBCUD4F_8|PDEN VSS BBCUD4F_5|Y BBCUD4F_9|PUEN VDD3V3 VDD3V3 BBCUD4F_2|A  ICF_2|PI comp_inp SCK gpio<9> ICFC_0|VDD3 BBC4F_3|A VDD1V8 BBCUD4F_14|PI BBCUD4F_0|EN  flash_io0 VDD1V8 comp_inp VDD1V8 VDD1V8 BBCUD4F_7|PI BBC4F_1|PI VDD3V3 BBCUD4F_0|PDEN  ICF_1|Y gpio<14> BBCUD4F_13|Y VDD1V8 BBCUD4F_1|PUEN BT4F_2|A BBCUD4F_13|PDEN VDD1V8  VDD3V3 VDD1V8 VDD3V3 BBCUD4F_10|A VDD1V8 gpio<2> BBCUD4F_14|PUEN VDD3V3 BBCUD4F_9|Y  VDD1V8 VDD3V3 VDD1V8 BT4F_2|EN BBCUD4F_6|A VDD1V8 irq VDD3V3 VDD1V8 BBCUD4F_10|PI  BBCUD4F_7|PDEN BBCUD4F_8|PUEN BBCUD4F_0|Y BBCUD4F_14|EN VDD3V3 BBCUD4F_3|PI BBC4F_1|EN  BBCUD4F_7|EN BBC4F_1|Y ICFC_0|PI VDD1V8 APR00DF_3|PAD VDD3V3 VDD3V3 BBCUD4F_14|A  VDD1V8 BT4FC_0|A VDD1V8 gpio<6> VDD3V3 BT4FC_0|EN VDD1V8 BBCUD4F_12|PDEN BBCUD4F_0|PUEN  VDD3V3 VDD3V3 VSS BBCUD4F_13|PUEN VDD1V8 axtoc02_3v3_0|CLK BBCUD4F_10|EN BBCUD4F_4|Y  BBCUD4F_3|EN VSS gpio<11> BBCUD4F_1|A VDD1V8 VDD3V3 SDI BBC4F_2|A BBCUD4F_6|PDEN  BBCUD4F_7|PUEN VDD3V3 VDD3V3 VDD3V3 ICF_1|PI XCLK ICF_0|Y BBCUD4F_12|Y adc0_in BT4F_1|A  ICFC_0|VDD3 BBCUD4F_13|PI axtoc02_3v3_0|EN BBCUD4F_8|Y VDD1V8 VDD1V8 w_n1073741817_n1073741817#  VDD3V3 BBCUD4F_6|PI BBC4F_0|PI BBCUD4F_5|A flash_io1 BBCUD4F_11|PDEN VDD3V3 BBCUD4F_12|PUEN  gpio<15> gpio<3> VDD1V8 VDD1V8 VDD1V8 BBC4F_0|Y BT4F_1|EN aregc01_3v3_1|EN VDD3V3  VDD1V8 VDD1V8 BBCUD4F_5|PDEN VDD3V3 VDD1V8 BBCUD4F_6|PUEN ICFC_2|Y BBCUD4F_13|A  BBCUD4F_13|EN VDD1V8 VDD3V3 BBCUD4F_2|PI SDO BBC4F_0|EN BBCUD4F_6|EN BBCUD4F_9|A  ser_tx VDD3V3 axtoc02_3v3_0|XI VDD1V8 APR00DF_4|PAD BBCUD4F_3|Y aregc01_3v3_0|ENB  gpio<7> BBCUD4F_0|A VDD1V8 VDD3V3 BBCUD4F_10|PDEN adc1_in VDD3V3 BBC4F_1|A BBCUD4F_11|PUEN  VDD3V3 VDD1V8 VDD1V8 BBCUD4F_2|EN VDD1V8 VDD1V8 VDD3V3 BBCUD4F_9|PI BBC4F_3|PI gpio<12>  VDD3V3 ICFC_0|VDD3 BBCUD4F_11|Y gpio<0> BT4F_0|A VDD1V8 VDD3V3 BBCUD4F_5|PUEN BBCUD4F_4|PDEN  BBCUD4F_7|Y VDD3V3 flash_csb BBCUD4F_4|A VDD3V3 ICF_0|PI VDD1V8 VSS BBCUD4F_12|PI  adc1_in BBCUD4F_5|PI VDD3V3 VDD1V8 VDD3V3 ICFC_2|PI BBC4F_3|EN BBCUD4F_9|EN VDD1V8  axtoc02_3v3_0|XO BBCUD4F_10|PUEN flash_io3 BBCUD4F_15|Y VDD3V3 VDD3V3 aregc01_3v3_0|OUT  BBCUD4F_12|A ICFC_1|Y VDD3V3 gpio<4> VDD3V3 VDD1V8 BT4F_0|EN aregc01_3v3_0|EN BBCUD4F_8|A  flash_clk ICFC_0|VDD3 VDD1V8 BBCUD4F_3|PDEN BBCUD4F_4|PUEN VDD1V8 BBCUD4F_12|EN  BBCUD4F_2|Y VDD3V3 BBCUD4F_1|PI BBC4F_3|Y flash_io0 VDD1V8 BBCUD4F_5|EN VDD3V3 BBC4F_0|A  flash_io1 VDD3V3 VDD3V3 comp_inn XI adc0_in flash_io2 gpio<8> aregc01_3v3_1|ENB  VDD1V8 VDD1V8 BBCUD4F_10|Y VDD1V8 VDD1V8 flash_io3 BBCUD4F_6|Y BBCUD4F_15|PI BBCUD4F_1|EN  VDD3V3 BBCUD4F_8|PI BBC4F_2|PI BBCUD4F_3|A ICFC_0|VDD3 VDD1V8 gpio<13> VDD1V8 VDD1V8  VDD1V8 BBCUD4F_3|PUEN BBCUD4F_2|PDEN gpio<1> BBCUD4F_15|PDEN VDD1V8 VDD3V3 aregc01_3v3_1|VIN3  VDD3V3 VDD1V8 CSB ICF_2|Y BBCUD4F_14|Y VDD3V3 VDD1V8 BBCUD4F_11|PI ICFC_0|Y flash_clk  BBCUD4F_11|A BBCUD4F_9|PDEN BBCUD4F_15|EN ICFC_0|VDD3 VDD1V8 VDD3V3 VSS BBCUD4F_4|PI  ser_rx BBCUD4F_8|EN BBC4F_2|EN VDD1V8 ICFC_1|PI APR00DF_2|PAD BBCUD4F_7|A VDD3V3  VDD1V8 VDD3V3 XO flash_io2 gpio<5> BBCUD4F_1|Y VDD3V3 VSS aregc01_3v3_1|OUT BBC4F_2|Y  VDD1V8 BBCUD4F_1|PDEN VDD3V3 VDD3V3 BBCUD4F_14|PDEN BBCUD4F_15|PUEN flash_csb BBCUD4F_2|PUEN  VDD3V3 aregc01_3v3_0|VIN3 BBCUD4F_11|EN BBCUD4F_15|A
XCORNERESDF_3 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER01F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER01F
XFILLER10F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER10F
XFILLER20F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XFILLER50F_2 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XVDDPADF_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 VDDPADF
XVDDORPADF_4 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_3 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XICF_2 ICF_2|PO ICF_2|PI ICF_2|Y XCLK VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XBT4F_1 BT4F_1|EN BT4F_1|A flash_clk VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XBT4F_2 BT4F_2|EN BT4F_2|A flash_csb VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XBBC4F_0 BBC4F_0|EN BBC4F_0|A BBC4F_0|Y BBC4F_0|PO BBC4F_0|PI flash_io0 VDD3V3 VSS  VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_1 BBC4F_1|EN BBC4F_1|A BBC4F_1|Y BBC4F_1|PO BBC4F_1|PI flash_io1 VDD3V3 VSS  VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_3 BBC4F_3|EN BBC4F_3|A BBC4F_3|Y BBC4F_3|PO BBC4F_3|PI flash_io2 VDD3V3 VSS  VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_2 BBC4F_2|EN BBC4F_2|A BBC4F_2|Y BBC4F_2|PO BBC4F_2|PI flash_io3 VDD3V3 VSS  VSS VDD3V3 VDD1V8 BBC4F
XFILLER40F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER40F
XPOWERCUTVDD3FC_1 VDD3V3 VDD3V3 VSS VSS POWERCUTVDD3FC
XVDDPADFC_0 VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 VDDPADFC
XBT4FC_0 BT4FC_0|EN BT4FC_0|A SDO VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 BT4FC
XICFC_2 ICFC_2|PO ICFC_2|PI ICFC_2|Y SCK VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 ICFC
XICFC_1 ICFC_1|PO ICFC_1|PI ICFC_1|Y CSB VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 ICFC
XFILLER20FC_0 VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 FILLER20FC
XICFC_0 ICFC_0|PO ICFC_0|PI ICFC_0|Y SDI VDD3V3 VDD3V3 VSS VSS ICFC_0|VDD3 ICFC
XPOWERCUTVDD3FC_0 VDD3V3 VDD3V3 VSS VSS POWERCUTVDD3FC
XFILLER20F_8 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XBBCUD4F_15 BBCUD4F_15|EN BBCUD4F_15|A BBCUD4F_15|Y BBCUD4F_15|PO BBCUD4F_15|PI BBCUD4F_15|PUEN  BBCUD4F_15|PDEN gpio<15> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XGNDORPADF_5 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER20F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_2 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER20F_7 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XICF_0 ICF_0|PO ICF_0|PI ICF_0|Y ser_rx VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XBT4F_0 BT4F_0|EN BT4F_0|A ser_tx VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XICF_1 ICF_1|PO ICF_1|PI ICF_1|Y irq VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XAPR00DF_6 comp_inp VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_5 comp_inn VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XFILLER50F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XGNDORPADF_0 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XVDDORPADF_0 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XVDDPADF_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 VDDPADF
XFILLER20F_6 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XGNDORPADF_2 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER50F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XGNDORPADF_6 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XVDDORPADF_2 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XFILLER01F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER01F
XBBCUD4F_14 BBCUD4F_14|EN BBCUD4F_14|A BBCUD4F_14|Y BBCUD4F_14|PO BBCUD4F_14|PI BBCUD4F_14|PUEN  BBCUD4F_14|PDEN gpio<14> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_13 BBCUD4F_13|EN BBCUD4F_13|A BBCUD4F_13|Y BBCUD4F_13|PO BBCUD4F_13|PI BBCUD4F_13|PUEN  BBCUD4F_13|PDEN gpio<13> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_12 BBCUD4F_12|EN BBCUD4F_12|A BBCUD4F_12|Y BBCUD4F_12|PO BBCUD4F_12|PI BBCUD4F_12|PUEN  BBCUD4F_12|PDEN gpio<12> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_11 BBCUD4F_11|EN BBCUD4F_11|A BBCUD4F_11|Y BBCUD4F_11|PO BBCUD4F_11|PI BBCUD4F_11|PUEN  BBCUD4F_11|PDEN gpio<11> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_10 BBCUD4F_10|EN BBCUD4F_10|A BBCUD4F_10|Y BBCUD4F_10|PO BBCUD4F_10|PI BBCUD4F_10|PUEN  BBCUD4F_10|PDEN gpio<10> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_9 BBCUD4F_9|EN BBCUD4F_9|A BBCUD4F_9|Y BBCUD4F_9|PO BBCUD4F_9|PI BBCUD4F_9|PUEN  BBCUD4F_9|PDEN gpio<9> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_8 BBCUD4F_8|EN BBCUD4F_8|A BBCUD4F_8|Y BBCUD4F_8|PO BBCUD4F_8|PI BBCUD4F_8|PUEN  BBCUD4F_8|PDEN gpio<8> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_7 BBCUD4F_7|EN BBCUD4F_7|A BBCUD4F_7|Y BBCUD4F_7|PO BBCUD4F_7|PI BBCUD4F_7|PUEN  BBCUD4F_7|PDEN gpio<7> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
Xaregc01_3v3_1 aregc01_3v3_1|OUT aregc01_3v3_1|EN aregc01_3v3_1|VIN3 aregc01_3v3_1|ENB  VDD1V8 VDD3V3 VSS VSS VDD3V3 aregc01_3v3
XBBCUD4F_6 BBCUD4F_6|EN BBCUD4F_6|A BBCUD4F_6|Y BBCUD4F_6|PO BBCUD4F_6|PI BBCUD4F_6|PUEN  BBCUD4F_6|PDEN gpio<6> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_5 BBCUD4F_5|EN BBCUD4F_5|A BBCUD4F_5|Y BBCUD4F_5|PO BBCUD4F_5|PI BBCUD4F_5|PUEN  BBCUD4F_5|PDEN gpio<5> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_4 BBCUD4F_4|EN BBCUD4F_4|A BBCUD4F_4|Y BBCUD4F_4|PO BBCUD4F_4|PI BBCUD4F_4|PUEN  BBCUD4F_4|PDEN gpio<4> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_3 BBCUD4F_3|EN BBCUD4F_3|A BBCUD4F_3|Y BBCUD4F_3|PO BBCUD4F_3|PI BBCUD4F_3|PUEN  BBCUD4F_3|PDEN gpio<3> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XFILLER20F_4 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_0 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER20F_2 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XAPR00DF_4 APR00DF_4|PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_3 APR00DF_3|PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_2 APR00DF_2|PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_1 adc1_in VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_0 adc0_in VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XVDDORPADF_1 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_1 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
Xaregc01_3v3_0 aregc01_3v3_0|OUT aregc01_3v3_0|EN aregc01_3v3_0|VIN3 aregc01_3v3_0|ENB  VDD1V8 VDD3V3 VSS VSS VDD3V3 aregc01_3v3
XFILLER20F_5 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XFILLER10F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER10F
XFILLER02F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER02F
XVDDORPADF_3 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_7 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER02F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER02F
Xaxtoc02_3v3_0 VSS VDD3V3 VSS VDD3V3 VDD1V8 axtoc02_3v3_0|XI axtoc02_3v3_0|XO axtoc02_3v3_0|CLK  axtoc02_3v3_0|EN axtoc02_3v3
XBBCUD4F_1 BBCUD4F_1|EN BBCUD4F_1|A BBCUD4F_1|Y BBCUD4F_1|PO BBCUD4F_1|PI BBCUD4F_1|PUEN  BBCUD4F_1|PDEN gpio<0> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_0 BBCUD4F_0|EN BBCUD4F_0|A BBCUD4F_0|Y BBCUD4F_0|PO BBCUD4F_0|PI BBCUD4F_0|PUEN  BBCUD4F_0|PDEN gpio<1> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_2 BBCUD4F_2|EN BBCUD4F_2|A BBCUD4F_2|Y BBCUD4F_2|PO BBCUD4F_2|PI BBCUD4F_2|PUEN  BBCUD4F_2|PDEN gpio<2> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XFILLER20F_3 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_1 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
C0 BBCUD4F_4|PI BBCUD4F_4|Y 0.01fF
C1 BBCUD4F_14|PI BBCUD4F_14|Y 0.01fF
C2 ICFC_0|PI ICFC_0|PO 0.04fF
C3 BT4FC_0|A BT4FC_0|EN 0.04fF
C4 axtoc02_3v3_0|m4_0_28769# axtoc02_3v3_0|m4_0_22024# 0.09fF
C5 BBCUD4F_13|A BBCUD4F_13|EN 0.04fF
C6 BBCUD4F_6|PI BBCUD4F_6|PO 0.04fF
C7 BBCUD4F_7|PDEN BBCUD4F_7|PUEN 0.04fF
C8 VDD3V3 axtoc02_3v3_0|m4_0_30653# 0.22fF
C9 BBCUD4F_7|A BBCUD4F_7|EN 0.04fF
C10 BBCUD4F_0|PI BBCUD4F_0|PO 0.04fF
C11 axtoc02_3v3_0|m4_0_31172# axtoc02_3v3_0|m4_0_30653# 0.26fF
C12 BBCUD4F_5|PI BBCUD4F_5|Y 0.01fF
C13 BBC4F_1|A BBC4F_1|EN 0.04fF
C14 BBC4F_3|A BBC4F_3|EN 0.04fF
C15 BBCUD4F_4|PO BBCUD4F_4|Y 0.04fF
C16 ICFC_0|PI ICFC_0|Y 0.01fF
C17 VDD3V3 axtoc02_3v3_0|m4_0_22024# 3.50fF
C18 BBCUD4F_6|PI BBCUD4F_6|Y 0.01fF
C19 axtoc02_3v3_0|m4_0_29333# axtoc02_3v3_0|m4_0_29057# 0.33fF
C20 axtoc02_3v3_0|m4_0_30133# axtoc02_3v3_0|m4_0_28769# 0.03fF
C21 axtoc02_3v3_0|m4_0_28769# VSS 0.11fF
C22 BBCUD4F_2|PI BBCUD4F_2|PO 0.04fF
C23 BBC4F_0|A BBC4F_0|EN 0.04fF
C24 BBCUD4F_15|PI BBCUD4F_15|Y 0.01fF
C25 BBCUD4F_5|PO BBCUD4F_5|Y 0.04fF
C26 VDD1V8 VSS 17.44fF
C27 ICF_0|PO ICF_0|Y 0.04fF
C28 BBCUD4F_12|PDEN BBCUD4F_12|PUEN 0.04fF
C29 ICF_2|PI ICF_2|PO 0.04fF
C30 BBCUD4F_8|PDEN BBCUD4F_8|PUEN 0.04fF
C31 BBCUD4F_11|PO BBCUD4F_11|Y 0.04fF
C32 BBCUD4F_12|PI BBCUD4F_12|PO 0.04fF
C33 BBCUD4F_14|PO BBCUD4F_14|Y 0.04fF
C34 BBCUD4F_8|A BBCUD4F_8|EN 0.04fF
C35 ICFC_0|PO ICFC_0|Y 0.04fF
C36 BBCUD4F_6|PO BBCUD4F_6|Y 0.04fF
C37 BBCUD4F_1|PDEN BBCUD4F_1|PUEN 0.04fF
C38 BBCUD4F_0|PI BBCUD4F_0|Y 0.01fF
C39 VDD3V3 VSS 260.23fF
C40 BBCUD4F_2|PI BBCUD4F_2|Y 0.01fF
C41 axtoc02_3v3_0|m4_0_31172# axtoc02_3v3_0|m4_0_30133# 0.05fF
C42 BBCUD4F_9|PDEN BBCUD4F_9|PUEN 0.04fF
C43 BBCUD4F_15|PO BBCUD4F_15|Y 0.04fF
C44 BBCUD4F_9|A BBCUD4F_9|EN 0.04fF
C45 ICF_2|PI ICF_2|Y 0.01fF
C46 BBCUD4F_12|PI BBCUD4F_12|Y 0.01fF
C47 BT4F_0|A BT4F_0|EN 0.04fF
C48 BT4F_2|A BT4F_2|EN 0.04fF
C49 BBCUD4F_11|A BBCUD4F_11|EN 0.04fF
C50 BBCUD4F_10|PDEN BBCUD4F_10|PUEN 0.04fF
C51 ICF_1|PI ICF_1|PO 0.04fF
C52 ICFC_0|VDD3 VSS 1.43fF
C53 BBCUD4F_14|A BBCUD4F_14|EN 0.04fF
C54 axtoc02_3v3_0|m4_0_29333# axtoc02_3v3_0|m4_0_28769# 0.08fF
C55 BBCUD4F_3|PDEN BBCUD4F_3|PUEN 0.04fF
C56 BBCUD4F_10|A BBCUD4F_10|EN 0.04fF
C57 BBCUD4F_0|PO BBCUD4F_0|Y 0.04fF
C58 BBCUD4F_2|PO BBCUD4F_2|Y 0.04fF
C59 BBCUD4F_1|PI BBCUD4F_1|PO 0.04fF
C60 BBCUD4F_3|A BBCUD4F_3|EN 0.04fF
C61 ICFC_2|PI ICFC_2|PO 0.04fF
C62 BT4F_1|A BT4F_1|EN 0.04fF
C63 BBCUD4F_15|A BBCUD4F_15|EN 0.04fF
C64 ICF_2|PO ICF_2|Y 0.04fF
C65 axtoc02_3v3_0|m4_0_29057# axtoc02_3v3_0|m4_0_28769# 0.33fF
C66 BBCUD4F_7|PI BBCUD4F_7|PO 0.04fF
C67 ICFC_2|PI ICFC_2|Y 0.01fF
C68 axtoc02_3v3_0|m4_0_30653# axtoc02_3v3_0|m4_0_30133# 0.26fF
C69 axtoc02_3v3_0|m4_0_31172# axtoc02_3v3_0|m4_0_29333# 0.03fF
C70 BBCUD4F_0|A BBCUD4F_0|EN 0.04fF
C71 BBCUD4F_15|A VSS 0.01fF
C72 ICFC_1|PI ICFC_1|PO 0.04fF
C73 BBCUD4F_12|PO BBCUD4F_12|Y 0.04fF
C74 BBCUD4F_4|PDEN BBCUD4F_4|PUEN 0.04fF
C75 ICF_1|PI ICF_1|Y 0.01fF
C76 BBCUD4F_4|A BBCUD4F_4|EN 0.04fF
C77 VDD3V3 axtoc02_3v3_0|m4_0_29057# 0.11fF
C78 BBCUD4F_7|PI BBCUD4F_7|Y 0.01fF
C79 ICFC_2|PO ICFC_2|Y 0.04fF
C80 BBC4F_0|PI BBC4F_0|PO 0.04fF
C81 BBCUD4F_1|PI BBCUD4F_1|Y 0.01fF
C82 axtoc02_3v3_0|XO XO 7.60fF
C83 axtoc02_3v3_0|XI XI 7.60fF
C84 BBCUD4F_5|PDEN BBCUD4F_5|PUEN 0.04fF
C85 BBCUD4F_5|A BBCUD4F_5|EN 0.04fF
C86 aregc01_3v3_1|ENB aregc01_3v3_1|VIN3 0.01fF
C87 BBC4F_2|PI BBC4F_2|PO 0.04fF
C88 ICFC_1|PI ICFC_1|Y 0.01fF
C89 BBCUD4F_13|PDEN BBCUD4F_13|PUEN 0.04fF
C90 BBCUD4F_8|PI BBCUD4F_8|PO 0.04fF
C91 BBCUD4F_12|A BBCUD4F_12|EN 0.04fF
C92 ICF_1|PO ICF_1|Y 0.04fF
C93 BBCUD4F_13|PI BBCUD4F_13|PO 0.04fF
C94 BBCUD4F_6|PDEN BBCUD4F_6|PUEN 0.04fF
C95 BBCUD4F_6|A BBCUD4F_6|EN 0.04fF
C96 BBCUD4F_7|PO BBCUD4F_7|Y 0.04fF
C97 BBC4F_0|PI BBC4F_0|Y 0.01fF
C98 BBCUD4F_1|PO BBCUD4F_1|Y 0.04fF
C99 axtoc02_3v3_0|m4_0_30653# axtoc02_3v3_0|m4_0_29333# 0.05fF
C100 axtoc02_3v3_0|m4_0_30133# VSS 0.22fF
C101 BBCUD4F_9|PI BBCUD4F_9|PO 0.04fF
C102 BBC4F_1|PI BBC4F_1|PO 0.04fF
C103 aregc01_3v3_0|ENB aregc01_3v3_0|VIN3 0.01fF
C104 aregc01_3v3_1|EN aregc01_3v3_1|VIN3 0.01fF
C105 BBC4F_3|PI BBC4F_3|PO 0.04fF
C106 ICFC_1|PO ICFC_1|Y 0.04fF
C107 aregc01_3v3_1|ENB aregc01_3v3_1|EN 0.06fF
C108 BBCUD4F_8|PI BBCUD4F_8|Y 0.01fF
C109 BBCUD4F_13|PI BBCUD4F_13|Y 0.01fF
C110 BBCUD4F_10|PI BBCUD4F_10|PO 0.04fF
C111 axtoc02_3v3_0|m4_0_29333# axtoc02_3v3_0|m4_0_22024# 0.03fF
C112 BBCUD4F_3|PI BBCUD4F_3|PO 0.04fF
C113 BBC4F_0|PO BBC4F_0|Y 0.04fF
C114 BBCUD4F_2|PDEN BBCUD4F_2|PUEN 0.04fF
C115 axtoc02_3v3_0|m4_0_30653# axtoc02_3v3_0|m4_0_29057# 0.02fF
C116 BBCUD4F_2|A BBCUD4F_2|EN 0.04fF
C117 BBCUD4F_1|A BBCUD4F_1|EN 0.04fF
C118 VDD1V8 VDD3V3 52.10fF
C119 BBCUD4F_9|PI BBCUD4F_9|Y 0.01fF
C120 VDD1V8 axtoc02_3v3_0|m4_0_31172# 0.37fF
C121 aregc01_3v3_0|EN aregc01_3v3_0|VIN3 0.01fF
C122 BBC4F_2|PI BBC4F_2|Y 0.01fF
C123 BBC4F_3|PI BBC4F_3|Y 0.01fF
C124 BBCUD4F_8|PO BBCUD4F_8|Y 0.04fF
C125 axtoc02_3v3_0|m4_0_29057# axtoc02_3v3_0|m4_0_22024# 0.05fF
C126 BBCUD4F_10|PI BBCUD4F_10|Y 0.01fF
C127 ICFC_0|VDD3 VDD1V8 0.67fF
C128 axtoc02_3v3_0|m4_0_0# VSS 3.72fF
C129 axtoc02_3v3_0|m4_0_30133# axtoc02_3v3_0|m4_0_29333# 0.26fF
C130 BBCUD4F_3|PI BBCUD4F_3|Y 0.01fF
C131 axtoc02_3v3_0|m4_0_29333# VSS 0.37fF
C132 BBCUD4F_15|PDEN BBCUD4F_15|PUEN 0.04fF
C133 BBCUD4F_9|PO BBCUD4F_9|Y 0.04fF
C134 BBC4F_1|PI BBC4F_1|Y 0.01fF
C135 BBC4F_2|PO BBC4F_2|Y 0.04fF
C136 ICF_0|PI ICF_0|PO 0.04fF
C137 BBCUD4F_11|PDEN BBCUD4F_11|PUEN 0.04fF
C138 aregc01_3v3_0|ENB aregc01_3v3_0|EN 0.06fF
C139 BBCUD4F_14|PDEN BBCUD4F_14|PUEN 0.04fF
C140 ICFC_0|VDD3 VDD3V3 4.25fF
C141 BBCUD4F_11|PI BBCUD4F_11|PO 0.04fF
C142 BBCUD4F_4|PI BBCUD4F_4|PO 0.04fF
C143 BBCUD4F_13|PO BBCUD4F_13|Y 0.04fF
C144 BBCUD4F_14|PI BBCUD4F_14|PO 0.04fF
C145 BBCUD4F_10|PO BBCUD4F_10|Y 0.04fF
C146 BBCUD4F_0|PDEN BBCUD4F_0|PUEN 0.04fF
C147 axtoc02_3v3_0|m4_0_30133# axtoc02_3v3_0|m4_0_29057# 0.03fF
C148 BBCUD4F_3|PO BBCUD4F_3|Y 0.04fF
C149 BBCUD4F_15|PI BBCUD4F_15|PO 0.04fF
C150 BBCUD4F_5|PI BBCUD4F_5|PO 0.04fF
C151 BBC4F_1|PO BBC4F_1|Y 0.04fF
C152 ICF_0|PI ICF_0|Y 0.01fF
C153 BBC4F_3|PO BBC4F_3|Y 0.04fF
C154 BBC4F_2|A BBC4F_2|EN 0.04fF
C155 BBCUD4F_11|PI BBCUD4F_11|Y 0.01fF
C156 XI w_n1073741817_n1073741817# -2.82fF
C157 XO w_n1073741817_n1073741817# -2.82fF
C158 gpio<2> w_n1073741817_n1073741817# -49.46fF
C159 gpio<1> w_n1073741817_n1073741817# 3.06fF
C160 gpio<0> w_n1073741817_n1073741817# 6.15fF
C161 VSS w_n1073741817_n1073741817# 32.97fF
C162 adc0_in w_n1073741817_n1073741817# 32.97fF
C163 adc1_in w_n1073741817_n1073741817# 32.97fF
C164 APR00DF_2|PAD w_n1073741817_n1073741817# 32.97fF
C165 APR00DF_3|PAD w_n1073741817_n1073741817# 32.97fF
C166 APR00DF_4|PAD w_n1073741817_n1073741817# 15.35fF
C167 gpio<3> w_n1073741817_n1073741817# 32.97fF
C168 gpio<4> w_n1073741817_n1073741817# 25.15fF
C169 gpio<5> w_n1073741817_n1073741817# 32.97fF
C170 gpio<6> w_n1073741817_n1073741817# 32.97fF
C171 VDD3V3 w_n1073741817_n1073741817# 32.97fF
C172 VDD1V8 w_n1073741817_n1073741817# 32.97fF
C173 gpio<7> w_n1073741817_n1073741817# 32.97fF
C174 gpio<8> w_n1073741817_n1073741817# 32.97fF
C175 gpio<9> w_n1073741817_n1073741817# 32.97fF
C176 gpio<10> w_n1073741817_n1073741817# 31.51fF
C177 gpio<11> w_n1073741817_n1073741817# 6.06fF
C178 gpio<12> w_n1073741817_n1073741817# 32.97fF
C179 gpio<13> w_n1073741817_n1073741817# 32.97fF
C180 gpio<14> w_n1073741817_n1073741817# 32.97fF
C181 comp_inn w_n1073741817_n1073741817# 32.97fF
C182 comp_inp w_n1073741817_n1073741817# 32.97fF
C183 irq w_n1073741817_n1073741817# 32.97fF
C184 ser_tx w_n1073741817_n1073741817# 32.97fF
C185 ser_rx w_n1073741817_n1073741817# 8.32fF
C186 gpio<15> w_n1073741817_n1073741817# 32.97fF
C187 SDI w_n1073741817_n1073741817# 18.78fF
C188 CSB w_n1073741817_n1073741817# 12.42fF
C189 SCK w_n1073741817_n1073741817# 32.97fF
C190 SDO w_n1073741817_n1073741817# 32.97fF
C191 flash_io3 w_n1073741817_n1073741817# 32.97fF
C192 flash_io2 w_n1073741817_n1073741817# 32.97fF
C193 flash_io1 w_n1073741817_n1073741817# 32.97fF
C194 flash_io0 w_n1073741817_n1073741817# 32.97fF
C195 flash_csb w_n1073741817_n1073741817# 32.97fF
C196 flash_clk w_n1073741817_n1073741817# 10.83fF
C197 XCLK w_n1073741817_n1073741817# 32.97fF
.ends

* Need include to schematic netlist for LOGIC0_3V

* Need include to schematic netlist for LOGIC1_3V

* Black-box entry replaced by path to RCX netlist
.include /home/wflisseg/design/ip/AMUX4_3V/11.0/spi-rcx/AMUX4_3V/AMUX4_3V__AMUX4_3V.spi

* Black-box entry replaced by path to schematic netlist
.include /home/wflisseg/design/ip/XSPRAM_1024X32_M8P/3.0/spi/XSPRAM_1024X32_M8P.spi

* Need include to schematic netlist for abgpc01_3v3
* Unknown black-box entry abgpc01_3v3
.subckt abgpc01_3v3 VDDA VSSA EN VBGVTN VBGP

* Need include to schematic netlist for acmpc01_3v3
* Unknown black-box entry acmpc01_3v3
.subckt acmpc01_3v3 IBN INP INN EN OUT VDDA VSSA

* Need include to schematic netlist for acsoc01_3v3
* Unknown black-box entry acsoc01_3v3
.subckt acsoc01_3v3 VDDA VSSA EN CS2_200N CS1_200N CS0_200N CS3_200N

* Need include to schematic netlist for arcoc01_3v3
* Unknown black-box entry arcoc01_3v3
.subckt arcoc01_3v3 EN CLK VDDA VSSA

* Need include to schematic netlist for aporc02_3v3
* Unknown black-box entry aporc02_3v3
.subckt aporc02_3v3 POR PORB VDDA VSSA

* Black-box entry replaced by path to RCX netlist
.include /home/wflisseg/design/ip/raven_spi/5.0/spi-rcx/raven_spi/raven_spi__raven_spi.spi

* Black-box entry replaced by path to RCX netlist
.include /home/wflisseg/design/ip/LS_3VX2/8.0/spi-rcx/LS_3VX2/LS_3VX2__LS_3VX2.spi

* Need include to schematic netlist for BU_3VX2

.subckt cmm5t_x3bss8 m4_2311_n4260# m4_6805_n4260# m4_24881_n4160# m4_29375_n4160#  m4_33869_n4160# w_n1073741817_n1073741817# m4_11399_n4160# m4_15893_n4160# m4_20387_n4160#  m4_n6677_n4260# m4_n2183_n4260# m4_n38135_n4260# m4_n33641_n4260# m4_n29147_n4260#  m4_6905_n4160# m4_n24653_n4260# m4_n20159_n4260# m4_n15665_n4260# m4_2411_n4160#  m4_n11171_n4260# m4_n6577_n4160# m4_n2083_n4160# m4_n38035_n4160# m4_n33541_n4160#  m4_n29047_n4160# m4_n24553_n4160# m4_n20059_n4160# m4_n15565_n4160# m4_n11071_n4160#  m4_24781_n4260# m4_29275_n4260# m4_33769_n4260# m4_11299_n4260# m4_15793_n4260#  m4_20287_n4260#
X0 m4_n38035_n4160# m4_n38135_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X1 m4_n33541_n4160# m4_n33641_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X2 m4_n29047_n4160# m4_n29147_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X3 m4_n24553_n4160# m4_n24653_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X4 m4_n20059_n4160# m4_n20159_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X5 m4_n15565_n4160# m4_n15665_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X6 m4_n11071_n4160# m4_n11171_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X7 m4_n6577_n4160# m4_n6677_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X8 m4_n2083_n4160# m4_n2183_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X9 m4_2411_n4160# m4_2311_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X10 m4_6905_n4160# m4_6805_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X11 m4_11399_n4160# m4_11299_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X12 m4_15893_n4160# m4_15793_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X13 m4_20387_n4160# m4_20287_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X14 m4_24881_n4160# m4_24781_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X15 m4_29375_n4160# m4_29275_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X16 m4_33869_n4160# m4_33769_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X17 m4_n38035_n4160# m4_n38135_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X18 m4_n33541_n4160# m4_n33641_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X19 m4_n29047_n4160# m4_n29147_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X20 m4_n24553_n4160# m4_n24653_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X21 m4_n20059_n4160# m4_n20159_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X22 m4_n15565_n4160# m4_n15665_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X23 m4_n11071_n4160# m4_n11171_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X24 m4_n6577_n4160# m4_n6677_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X25 m4_n2083_n4160# m4_n2183_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X26 m4_2411_n4160# m4_2311_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X27 m4_6905_n4160# m4_6805_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X28 m4_11399_n4160# m4_11299_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X29 m4_15893_n4160# m4_15793_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X30 m4_20387_n4160# m4_20287_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X31 m4_24881_n4160# m4_24781_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X32 m4_29375_n4160# m4_29275_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X33 m4_33869_n4160# m4_33769_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
C0 m4_n24653_n4260# m4_n20159_n4260# 6.69fF
C1 m4_n33641_n4260# m4_n29047_n4160# 3.54fF
C2 m4_n29147_n4260# m4_n24653_n4260# 6.69fF
C3 m4_2411_n4160# m4_6905_n4160# 1.65fF
C4 m4_n2183_n4260# m4_n2083_n4160# 5.16fF
C5 m4_20287_n4260# m4_24881_n4160# 3.54fF
C6 m4_11299_n4260# m4_11399_n4160# 5.16fF
C7 m4_n24653_n4260# m4_n20059_n4160# 3.54fF
C8 m4_n15665_n4260# m4_n15565_n4160# 5.16fF
C9 m4_33769_n4260# m4_33869_n4160# 5.16fF
C10 m4_24781_n4260# m4_29275_n4260# 6.69fF
C11 m4_n38135_n4260# m4_n38035_n4160# 5.16fF
C12 m4_11299_n4260# m4_15793_n4260# 6.69fF
C13 m4_n20159_n4260# m4_n15665_n4260# 6.69fF
C14 m4_n15665_n4260# m4_n11171_n4260# 6.69fF
C15 m4_6805_n4260# m4_6905_n4160# 5.16fF
C16 m4_n2183_n4260# m4_2311_n4260# 6.69fF
C17 m4_24781_n4260# m4_29375_n4160# 3.54fF
C18 m4_n20159_n4260# m4_n15565_n4160# 3.54fF
C19 m4_n15665_n4260# m4_n11071_n4160# 3.54fF
C20 m4_n33541_n4160# m4_n29047_n4160# 1.65fF
C21 m4_n29147_n4260# m4_n24553_n4160# 3.54fF
C22 m4_n2183_n4260# m4_2411_n4160# 3.54fF
C23 m4_n38135_n4260# m4_n33641_n4260# 6.69fF
C24 m4_24881_n4160# m4_29375_n4160# 1.65fF
C25 m4_11299_n4260# m4_15893_n4160# 3.54fF
C26 m4_n24553_n4160# m4_n20059_n4160# 1.65fF
C27 m4_n6677_n4260# m4_n2183_n4260# 6.69fF
C28 m4_n20059_n4160# m4_n15565_n4160# 1.65fF
C29 m4_15793_n4260# m4_20387_n4160# 3.54fF
C30 m4_n15565_n4160# m4_n11071_n4160# 1.65fF
C31 m4_n2083_n4160# m4_2411_n4160# 1.65fF
C32 m4_n20159_n4260# m4_n20059_n4160# 5.16fF
C33 m4_n6677_n4260# m4_n2083_n4160# 3.54fF
C34 m4_6805_n4260# m4_11299_n4260# 6.69fF
C35 m4_n11171_n4260# m4_n11071_n4160# 5.16fF
C36 m4_n29147_n4260# m4_n33641_n4260# 6.69fF
C37 m4_29275_n4260# m4_29375_n4160# 5.16fF
C38 m4_11399_n4160# m4_15893_n4160# 1.65fF
C39 m4_n6577_n4160# m4_n2083_n4160# 1.65fF
C40 m4_15893_n4160# m4_20387_n4160# 1.65fF
C41 m4_n11171_n4260# m4_n6677_n4260# 6.69fF
C42 m4_n38135_n4260# m4_n33541_n4160# 3.54fF
C43 m4_2311_n4260# m4_2411_n4160# 5.16fF
C44 m4_15793_n4260# m4_15893_n4160# 5.16fF
C45 m4_20287_n4260# m4_20387_n4160# 5.16fF
C46 m4_20387_n4160# m4_24881_n4160# 1.65fF
C47 m4_6805_n4260# m4_11399_n4160# 3.54fF
C48 m4_n11171_n4260# m4_n6577_n4160# 3.54fF
C49 m4_n38035_n4160# m4_n33541_n4160# 1.65fF
C50 m4_29275_n4260# m4_33769_n4260# 6.69fF
C51 m4_15793_n4260# m4_20287_n4260# 6.69fF
C52 m4_n29047_n4160# m4_n24553_n4160# 1.65fF
C53 m4_6905_n4160# m4_11399_n4160# 1.65fF
C54 m4_n11071_n4160# m4_n6577_n4160# 1.65fF
C55 m4_2311_n4260# m4_6805_n4260# 6.69fF
C56 m4_29275_n4260# m4_33869_n4160# 3.54fF
C57 m4_n24653_n4260# m4_n24553_n4160# 5.16fF
C58 m4_n6677_n4260# m4_n6577_n4160# 5.16fF
C59 m4_n33641_n4260# m4_n33541_n4160# 5.16fF
C60 m4_n29147_n4260# m4_n29047_n4160# 5.16fF
C61 m4_2311_n4260# m4_6905_n4160# 3.54fF
C62 m4_29375_n4160# m4_33869_n4160# 1.65fF
C63 m4_20287_n4260# m4_24781_n4260# 6.69fF
C64 m4_24781_n4260# m4_24881_n4160# 5.16fF
C65 m4_33869_n4160# w_n1073741817_n1073741817# 4.82fF
C66 m4_33769_n4260# w_n1073741817_n1073741817# 1.79fF
C67 m4_29375_n4160# w_n1073741817_n1073741817# 4.82fF
C68 m4_29275_n4260# w_n1073741817_n1073741817# 1.79fF
C69 m4_24881_n4160# w_n1073741817_n1073741817# 4.82fF
C70 m4_24781_n4260# w_n1073741817_n1073741817# 1.79fF
C71 m4_20387_n4160# w_n1073741817_n1073741817# 4.82fF
C72 m4_20287_n4260# w_n1073741817_n1073741817# 1.79fF
C73 m4_15893_n4160# w_n1073741817_n1073741817# 4.82fF
C74 m4_15793_n4260# w_n1073741817_n1073741817# 1.79fF
C75 m4_11399_n4160# w_n1073741817_n1073741817# 4.82fF
C76 m4_11299_n4260# w_n1073741817_n1073741817# 1.79fF
C77 m4_6905_n4160# w_n1073741817_n1073741817# 4.82fF
C78 m4_6805_n4260# w_n1073741817_n1073741817# 1.79fF
C79 m4_2411_n4160# w_n1073741817_n1073741817# 4.82fF
C80 m4_2311_n4260# w_n1073741817_n1073741817# 1.79fF
C81 m4_n2083_n4160# w_n1073741817_n1073741817# 4.82fF
C82 m4_n2183_n4260# w_n1073741817_n1073741817# 1.79fF
C83 m4_n6577_n4160# w_n1073741817_n1073741817# 4.82fF
C84 m4_n6677_n4260# w_n1073741817_n1073741817# 1.79fF
C85 m4_n11071_n4160# w_n1073741817_n1073741817# 4.82fF
C86 m4_n11171_n4260# w_n1073741817_n1073741817# 1.79fF
C87 m4_n15565_n4160# w_n1073741817_n1073741817# 4.82fF
C88 m4_n15665_n4260# w_n1073741817_n1073741817# 1.79fF
C89 m4_n20059_n4160# w_n1073741817_n1073741817# 4.82fF
C90 m4_n20159_n4260# w_n1073741817_n1073741817# 1.79fF
C91 m4_n24553_n4160# w_n1073741817_n1073741817# 4.82fF
C92 m4_n24653_n4260# w_n1073741817_n1073741817# 1.79fF
C93 m4_n29047_n4160# w_n1073741817_n1073741817# 4.82fF
C94 m4_n29147_n4260# w_n1073741817_n1073741817# 1.79fF
C95 m4_n33541_n4160# w_n1073741817_n1073741817# 4.82fF
C96 m4_n33641_n4260# w_n1073741817_n1073741817# 1.79fF
C97 m4_n38035_n4160# w_n1073741817_n1073741817# 4.82fF
C98 m4_n38135_n4260# w_n1073741817_n1073741817# 1.79fF
.ends

* Need include to schematic netlist for atmpc01_3v3
* Unknown black-box entry atmpc01_3v3
.subckt atmpc01_3v3 OVT EN VSSA VDDA

* Need include to schematic netlist for aopac01_3v3
* Unknown black-box entry aopac01_3v3
.subckt aopac01_3v3 EN INP INN OUT IB VDDA VSSA

* Need include to schematic netlist for acsoc02_3v3
* Unknown black-box entry acsoc02_3v3
.subckt acsoc02_3v3 CS_2U CS_4U EN CS_1U CS_8U VSSA VDDA

* Black-box entry replaced by path to RCX netlist
.include /home/wflisseg/design/ip/AMUX2_3V/10.0/spi-rcx/AMUX2_3V/AMUX2_3V__AMUX2_3V.spi

* Need include to schematic netlist for adacc01_3v3
* Unknown black-box entry adacc01_3v3
.subckt adacc01_3v3 OUT VSSA VDDA D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0>  EN VSS VREFH VREFL VDD

* Black-box entry replaced by path to RCX netlist
.include /home/wflisseg/design/ip/raven_soc/11.0/spi-rcx/raven_soc/raven_soc__raven_soc.spi

* Need include to schematic netlist for aadcc01_3v3
* Unknown black-box entry aadcc01_3v3
.subckt aadcc01_3v3 VDD EOC EN START CLK D<0> D<1> D<2> D<3> D<4> D<5> D<6> D<7> D<8>  D<9> VIN VREFH VREFL VSSA VDDA VSS

* Need include to schematic netlist for IN_3VX2

* Need include to schematic netlist for apllc03_1v8
* Unknown black-box entry apllc03_1v8
.subckt apllc03_1v8 REF B_VCO B_CP VDDD VSSD B<3> B<2> B<1> B<0> VCO_IN CLK VSSA VDDA  EN_CP EN_VCO

* Need include to schematic netlist for acsoc04_1v8
* Unknown black-box entry acsoc04_1v8
.subckt acsoc04_1v8 CS1_2u EN VDDA VSSA CS0_1u CS2_4u CS3_8u

.subckt raven VDD3V3 vdd VSS XCLK SDI SDO CSB SCK ser_tx ser_rx irq gpio[15] gpio[14]  gpio[13] gpio[12] gpio[11] gpio[10] gpio[9] gpio[8] gpio[7] gpio[6] gpio[5] gpio[4]  gpio[3] gpio[2] gpio[1] gpio[0] flash_csb flash_clk flash_io0 flash_io1 flash_io2  flash_io3 adc_high adc_low adc0_in adc1_in analog_out comp_inp comp_inn XI XO adc0_data<5>
Xraven_padframe_0 raven_padframe_0|ICF_1|VDDR VDD LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<4>  gpio[10] VDD VDD3V3 XCLK comp_inn raven_soc_0|gpio_pulldown<8> VSS raven_soc_0|gpio_in<5>  raven_soc_0|gpio_pullup<9> raven_padframe_0|BBCUD4F_2|VDDR raven_padframe_0|BBCUD4F_15|VDDR  raven_soc_0|gpio_out<2> LOGIC0_3V_4|Q comp_inp SCK gpio[9] raven_padframe_0|FILLER20FC_0|VDD3  raven_soc_0|flash_io2_do VDD LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<1> flash_io0  VDD comp_inp VDD VDD LOGIC0_3V_4|Q LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_9|VDDR  raven_soc_0|gpio_pulldown<1> raven_soc_0|irq_pin gpio[14] raven_soc_0|gpio_in<13>  VDD raven_soc_0|gpio_pullup<0> raven_soc_0|flash_csb raven_soc_0|gpio_pulldown<13>  VDD raven_padframe_0|BBC4F_3|VDDR VDD raven_padframe_0|APR00DF_0|VDDR raven_soc_0|gpio_out<10>  vdd gpio[2] raven_soc_0|gpio_pullup<14> raven_padframe_0|ICF_0|VDDR raven_soc_0|gpio_in<9>  VDD VDD3V3 VDD LOGIC0_3V_4|Q raven_soc_0|gpio_out<6> VDD irq raven_padframe_0|FILLER40F_0|VDDR  VDD LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<1>  raven_soc_0|gpio_outenb<14> raven_padframe_0|BBCUD4F_14|VDDR LOGIC0_3V_4|Q raven_soc_0|flash_io1_oeb  raven_soc_0|gpio_outenb<7> raven_soc_0|flash_io1_di LOGIC0_3V_4|Q VDD adc_high raven_padframe_0|GNDORPADF_3|VDDR  raven_padframe_0|VDDPADFC_0|VDDR raven_soc_0|gpio_out<14> VDD raven_spi_0|SDO VDD  gpio[6] raven_padframe_0|BBCUD4F_8|VDDR raven_spi_0|sdo_enb VDD raven_soc_0|gpio_pulldown<12>  raven_soc_0|gpio_pullup<1> raven_padframe_0|BBC4F_2|VDDR raven_padframe_0|VDDPADF_1|VDDR  gnd raven_soc_0|gpio_pullup<13> VDD BU_3VX2_72|A raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<4>  raven_soc_0|gpio_outenb<3> gnd gpio[11] raven_soc_0|gpio_out<0> VDD raven_padframe_0|FILLER20F_5|VDDR  SDI raven_soc_0|flash_io3_do raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pullup<7>  raven_padframe_0|BBCUD4F_13|VDDR raven_padframe_0|BBCUD4F_0|VDDR VDD3V3 LOGIC0_3V_4|Q  XCLK raven_soc_0|ser_rx raven_soc_0|gpio_in<12> AMUX4_3V_0|AIN1 raven_soc_0|flash_clk  VDD3V3 LOGIC0_3V_4|Q BU_3VX2_31|A raven_soc_0|gpio_in<8> VDD VDD gnd raven_padframe_0|BBCUD4F_7|VDDR  LOGIC0_3V_4|Q LOGIC0_3V_4|Q raven_soc_0|gpio_out<5> flash_io1 raven_soc_0|gpio_pulldown<11>  raven_padframe_0|BBC4F_1|VDDR raven_soc_0|gpio_pullup<12> gpio[15] gpio[3] VDD VDD  VDD raven_soc_0|flash_io0_di LOGIC0_3V_4|Q IN_3VX2_1|A raven_padframe_0|ICFC_2|VDDR  VDD VDD raven_soc_0|gpio_pulldown<5> raven_padframe_0|FILLER02F_1|VDDR VDD raven_soc_0|gpio_pullup<6>  BU_3VX2_33|A raven_soc_0|gpio_out<13> raven_soc_0|gpio_outenb<13> VDD raven_padframe_0|BBCUD4F_12|VDDR  LOGIC0_3V_4|Q SDO raven_soc_0|flash_io0_oeb raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<9>  ser_tx raven_padframe_0|BT4F_2|VDDR raven_padframe_0|axtoc02_3v3_0|XI VDD analog_out  raven_soc_0|gpio_in<3> IN_3VX2_1|Q gpio[7] raven_soc_0|gpio_out<1> VDD raven_padframe_0|BBCUD4F_6|VDDR  raven_soc_0|gpio_pulldown<10> adc1_in raven_padframe_0|BBC4F_0|VDDR raven_soc_0|flash_io1_do  raven_soc_0|gpio_pullup<11> raven_padframe_0|POWERCUTVDD3FC_1|VDDR VDD VDD raven_soc_0|gpio_outenb<2>  VDD VDD raven_padframe_0|FILLER20F_3|VDDR LOGIC0_3V_4|Q LOGIC0_3V_4|Q gpio[12] raven_padframe_0|ICFC_1|VDDR  raven_padframe_0|ICFC_2|VDD3 raven_soc_0|gpio_in<11> gpio[0] raven_soc_0|ser_tx  VDD raven_padframe_0|FILLER02F_0|VDDR raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_pulldown<4>  raven_soc_0|gpio_in<7> raven_padframe_0|BBCUD4F_11|VDDR flash_csb raven_soc_0|gpio_out<4>  raven_padframe_0|BT4F_1|VDDR LOGIC0_3V_4|Q VDD gnd LOGIC0_3V_4|Q AMUX4_3V_1|AIN1  LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_5|VDDR VDD VDD3V3 LOGIC0_3V_4|Q raven_soc_0|flash_io2_oeb  raven_soc_0|gpio_outenb<9> VDD raven_padframe_0|axtoc02_3v3_0|XO raven_soc_0|gpio_pullup<10>  flash_io3 raven_soc_0|gpio_in<15> raven_padframe_0|POWERCUTVDD3FC_0|VDDR VDD3V3  vdd raven_soc_0|gpio_out<12> raven_spi_0|CSB raven_padframe_0|GNDORPADF_7|VDDR gpio[4]  raven_padframe_0|ICFC_0|VDDR VDD LOGIC0_3V_4|Q IN_3VX2_1|A raven_soc_0|gpio_out<8>  flash_clk raven_padframe_0|ICFC_1|VDD3 VDD raven_soc_0|gpio_pulldown<3> raven_soc_0|gpio_pullup<4>  VDD raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<2> raven_padframe_0|BBCUD4F_10|VDDR  LOGIC0_3V_4|Q raven_soc_0|flash_io2_di flash_io0 vdd raven_soc_0|gpio_outenb<5>  raven_padframe_0|BT4F_0|VDDR raven_soc_0|flash_io0_do flash_io1 raven_padframe_0|BT4FC_0|VDDR  raven_padframe_0|BBCUD4F_4|VDDR AMUX4_3V_4|AIN1 XI adc0_in flash_io2 gpio[8] IN_3VX2_1|Q  VDD VDD raven_soc_0|gpio_in<10> VDD VDD flash_io3 raven_soc_0|gpio_in<6> LOGIC0_3V_4|Q  raven_soc_0|gpio_outenb<0> raven_padframe_0|FILLER20F_1|VDDR LOGIC0_3V_4|Q LOGIC0_3V_4|Q  raven_soc_0|gpio_out<3> raven_padframe_0|ICFC_0|VDD3 VDD gpio[13] VDD VDD vdd raven_soc_0|gpio_pullup<3>  raven_soc_0|gpio_pulldown<2> gpio[1] raven_soc_0|gpio_pulldown<15> VDD raven_padframe_0|FILLER10F_0|VDDR  VDD3V3 raven_padframe_0|ICF_2|VDDR VDD CSB raven_soc_0|ext_clk raven_soc_0|gpio_in<14>  raven_padframe_0|FILLER20F_8|VDDR VDD LOGIC0_3V_4|Q raven_spi_0|SDI flash_clk raven_soc_0|gpio_out<11>  raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<15> raven_padframe_0|BT4FC_0|VDD3  VDD raven_padframe_0|BBCUD4F_3|VDDR gnd LOGIC0_3V_4|Q ser_rx raven_soc_0|gpio_outenb<8>  raven_soc_0|flash_io3_oeb VDD LOGIC0_3V_4|Q adc_low raven_soc_0|gpio_out<7> raven_padframe_0|FILLER20FC_0|VDDR  VDD raven_padframe_0|GNDORPADF_5|VDDR XO flash_io2 gpio[5] raven_soc_0|gpio_in<0>  raven_padframe_0|FILLER20F_0|VDDR gnd vdd raven_soc_0|flash_io3_di VDD raven_soc_0|gpio_pulldown<0>  raven_padframe_0|APR00DF_1|VDDR VDD3V3 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<15>  flash_csb raven_soc_0|gpio_pullup<2> raven_padframe_0|FILLER50F_2|VDDR VDD3V3 raven_soc_0|gpio_outenb<11>  raven_soc_0|gpio_out<15> raven_padframe
XLOGIC0_3V_4 LOGIC0_3V_4|Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_3 LOGIC0_3V_3|Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_2 LOGIC0_3V_2|Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_1 LOGIC0_3V_1|Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_0 LOGIC0_3V_0|Q gnd VDD3V3 LOGIC0_3V
XLOGIC1_3V_3 LOGIC1_3V_3|Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_2 LOGIC1_3V_2|Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_1 LOGIC1_3V_1|Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_0 LOGIC1_3V_0|Q gnd VDD3V3 LOGIC1_3V
XAMUX4_3V_3 comp_inp AMUX4_3V_4|AIN2 AMUX4_3V_4|AIN3 vdd AMUX4_3V_3|AOUT AMUX4_3V_3|SEL[1] AMUX4_3V_3|SEL[0] vdd VDD3V3 gnd AMUX4_3V__AMUX4_3V 
XAMUX4_3V_4 AMUX4_3V_4|AIN1 AMUX4_3V_4|AIN2 AMUX4_3V_4|AIN3 vdd AMUX4_3V_4|AOUT AMUX4_3V_4|SEL[1] AMUX4_3V_4|SEL[0] vdd VDD3V3 gnd AMUX4_3V__AMUX4_3V 
XXSPRAM_1024X32_M8P_0 raven_soc_0|ram_addr<0> raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<2>  raven_soc_0|ram_addr<3> raven_soc_0|ram_addr<4> raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<6>  raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<9> BU_3VX2_0|Q  apllc03_1v8_0|CLK raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<11>  raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<15>  raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<19>  raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<22>  raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<26>  raven_soc_0|ram_wdata<27> raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<29> raven_soc_0|ram_wdata<2>  raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<31> raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<4>  raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<8>  raven_soc_0|ram_wdata<9> BU_3VX2_0|Q raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<10>  raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<13> raven_soc_0|ram_rdata<14>  raven_soc_0|ram_rdata<15> raven_soc_0|ram_rdata<16> raven_soc_0|ram_rdata<17> raven_soc_0|ram_rdata<18>  raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<1> raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<21>  raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<25>  raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<29>  raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<3>  raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<7>  raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<9> XSPRAM_1024X32_M8P_0|RDY vdd gnd  raven_soc_0|ram_wenb XSPRAM_1024X32_M8P
Xabgpc01_3v3_0 VDD3V3 gnd LS_3VX2_18|Q abgpc01_3v3_0|VBGVTN AMUX4_3V_4|AIN3 abgpc01_3v3
Xacmpc01_3v3_0 acmpc01_3v3_0|IBN AMUX4_3V_3|AOUT AMUX4_3V_4|AOUT LS_3VX2_23|Q BU_3VX2_32|A  VDD3V3 gnd acmpc01_3v3
Xacsoc01_3v3_0 VDD3V3 gnd LS_3VX2_23|Q acsoc01_3v3_0|CS2_200N acmpc01_3v3_0|IBN acmpc01_3v3_0|IBN  acsoc01_3v3_0|CS3_200N acsoc01_3v3
Xarcoc01_3v3_0 LS_3VX2_2|Q BU_3VX2_1|A VDD3V3 gnd arcoc01_3v3
Xaporc02_3v3_0 BU_3VX2_0|A aporc02_3v3_0|PORB VDD3V3 gnd aporc02_3v3
Xraven_spi_0 VDD3V3 gnd BU_3VX2_0|A BU_3VX2_33|A raven_spi_0|SDI raven_spi_0|CSB LS_3VX2_3|Q LOGIC0_3V_0|Q LOGIC0_3V_1|Q LOGIC0_3V_2|Q LOGIC0_3V_3|Q raven_spi_0|SDO raven_spi_0|sdo_enb BU_3VX2_31|A IN_3VX2_1|A BU_3VX2_28|A BU_3VX2_29|A BU_3VX2_27|A BU_3VX2_26|A BU_3VX2_25|A BU_3VX2_24|A BU_3VX2_23|A BU_3VX2_40|A BU_3VX2_71|A BU_3VX2_63|A BU_3VX2_22|A BU_3VX2_21|A BU_3VX2_20|A BU_3VX2_19|A BU_3VX2_18|A BU_3VX2_17|A BU_3VX2_16|A BU_3VX2_15|A BU_3VX2_14|A BU_3VX2_13|A BU_3VX2_12|A BU_3VX2_11|A BU_3VX2_10|A BU_3VX2_9|A BU_3VX2_8|A BU_3VX2_7|A BU_3VX2_6|A BU_3VX2_5|A BU_3VX2_4|A BU_3VX2_3|A BU_3VX2_2|A BU_3VX2_37|A BU_3VX2_38|A BU_3VX2_35|A raven_spi__raven_spi 
XLS_3VX2_18 LS_3VX2_18|A LS_3VX2_18|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_23 LS_3VX2_23|A LS_3VX2_23|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_2 LS_3VX2_2|A LS_3VX2_2|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XBU_3VX2_70 BU_3VX2_70|A BU_3VX2_70|Q gnd vdd BU_3VX2
XBU_3VX2_69 BU_3VX2_69|A BU_3VX2_69|Q gnd vdd BU_3VX2
XBU_3VX2_68 BU_3VX2_68|A BU_3VX2_68|Q gnd vdd BU_3VX2
XBU_3VX2_67 BU_3VX2_67|A BU_3VX2_67|Q gnd vdd BU_3VX2
XBU_3VX2_66 BU_3VX2_66|A BU_3VX2_66|Q gnd vdd BU_3VX2
XBU_3VX2_65 BU_3VX2_65|A BU_3VX2_65|Q gnd vdd BU_3VX2
XBU_3VX2_64 BU_3VX2_64|A BU_3VX2_64|Q gnd vdd BU_3VX2
XBU_3VX2_36 BU_3VX2_36|A BU_3VX2_36|Q gnd vdd BU_3VX2
XBU_3VX2_1 BU_3VX2_1|A BU_3VX2_1|Q gnd vdd BU_3VX2
XBU_3VX2_33 BU_3VX2_33|A BU_3VX2_33|Q gnd vdd BU_3VX2
XBU_3VX2_32 BU_3VX2_32|A BU_3VX2_32|Q gnd vdd BU_3VX2
XLOGIC0_3V_12 BU_3VX2_70|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_11 BU_3VX2_69|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_10 BU_3VX2_68|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_9 BU_3VX2_67|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_8 BU_3VX2_66|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_7 BU_3VX2_65|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_6 BU_3VX2_64|A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_5 BU_3VX2_36|A gnd VDD3V3 LOGIC0_3V
XBU_3VX2_0 BU_3VX2_0|A BU_3VX2_0|Q gnd vdd BU_3VX2
XBU_3VX2_31 BU_3VX2_31|A BU_3VX2_31|Q gnd vdd BU_3VX2
XBU_3VX2_30 IN_3VX2_1|A BU_3VX2_30|Q gnd vdd BU_3VX2
XBU_3VX2_29 BU_3VX2_29|A BU_3VX2_29|Q gnd vdd BU_3VX2
XBU_3VX2_28 BU_3VX2_28|A BU_3VX2_28|Q gnd vdd BU_3VX2
XBU_3VX2_27 BU_3VX2_27|A BU_3VX2_27|Q gnd vdd BU_3VX2
XBU_3VX2_26 BU_3VX2_26|A BU_3VX2_26|Q gnd vdd BU_3VX2
XBU_3VX2_25 BU_3VX2_25|A BU_3VX2_25|Q gnd vdd BU_3VX2
XBU_3VX2_24 BU_3VX2_24|A BU_3VX2_24|Q gnd vdd BU_3VX2
XBU_3VX2_23 BU_3VX2_23|A BU_3VX2_23|Q gnd vdd BU_3VX2
XBU_3VX2_22 BU_3VX2_22|A BU_3VX2_22|Q gnd vdd BU_3VX2
XBU_3VX2_21 BU_3VX2_21|A BU_3VX2_21|Q gnd vdd BU_3VX2
XBU_3VX2_20 BU_3VX2_20|A BU_3VX2_20|Q gnd vdd BU_3VX2
XBU_3VX2_19 BU_3VX2_19|A BU_3VX2_19|Q gnd vdd BU_3VX2
XBU_3VX2_18 BU_3VX2_18|A BU_3VX2_18|Q gnd vdd BU_3VX2
XBU_3VX2_17 BU_3VX2_17|A BU_3VX2_17|Q gnd vdd BU_3VX2
XBU_3VX2_16 BU_3VX2_16|A BU_3VX2_16|Q gnd vdd BU_3VX2
XBU_3VX2_15 BU_3VX2_15|A BU_3VX2_15|Q gnd vdd BU_3VX2
XBU_3VX2_14 BU_3VX2_14|A BU_3VX2_14|Q gnd vdd BU_3VX2
XBU_3VX2_13 BU_3VX2_13|A BU_3VX2_13|Q gnd vdd BU_3VX2
XBU_3VX2_12 BU_3VX2_12|A BU_3VX2_12|Q gnd vdd BU_3VX2
XBU_3VX2_11 BU_3VX2_11|A BU_3VX2_11|Q gnd vdd BU_3VX2
XBU_3VX2_10 BU_3VX2_10|A BU_3VX2_10|Q gnd vdd BU_3VX2
XBU_3VX2_9 BU_3VX2_9|A BU_3VX2_9|Q gnd vdd BU_3VX2
XBU_3VX2_8 BU_3VX2_8|A BU_3VX2_8|Q gnd vdd BU_3VX2
XBU_3VX2_7 BU_3VX2_7|A BU_3VX2_7|Q gnd vdd BU_3VX2
XBU_3VX2_6 BU_3VX2_6|A BU_3VX2_6|Q gnd vdd BU_3VX2
XBU_3VX2_5 BU_3VX2_5|A BU_3VX2_5|Q gnd vdd BU_3VX2
XBU_3VX2_4 BU_3VX2_4|A BU_3VX2_4|Q gnd vdd BU_3VX2
XBU_3VX2_3 BU_3VX2_3|A BU_3VX2_3|Q gnd vdd BU_3VX2
XBU_3VX2_2 BU_3VX2_2|A BU_3VX2_2|Q gnd vdd BU_3VX2
XBU_3VX2_37 BU_3VX2_37|A BU_3VX2_37|Q gnd vdd BU_3VX2
XBU_3VX2_38 BU_3VX2_38|A BU_3VX2_38|Q gnd vdd BU_3VX2
XBU_3VX2_35 BU_3VX2_35|A BU_3VX2_35|Q gnd vdd BU_3VX2
XBU_3VX2_40 BU_3VX2_40|A BU_3VX2_40|Q gnd vdd BU_3VX2
XBU_3VX2_63 BU_3VX2_63|A BU_3VX2_63|Q gnd vdd BU_3VX2
XBU_3VX2_71 BU_3VX2_71|A BU_3VX2_71|Q gnd vdd BU_3VX2
XLS_3VX2_3 LS_3VX2_3|A LS_3VX2_3|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
Xcmm5t_x3bss8_0 gnd gnd VDD3V3 VDD3V3 VDD3V3 gnd VDD3V3 VDD3V3 VDD3V3 gnd gnd gnd  gnd gnd VDD3V3 gnd gnd gnd VDD3V3 gnd VDD3V3 VDD3V3 VDD3V3 VDD3V3 VDD3V3 VDD3V3  VDD3V3 VDD3V3 VDD3V3 gnd gnd gnd gnd gnd gnd cmm5t_x3bss8
Xatmpc01_3v3_0 BU_3VX2_73|A LS_3VX2_24|Q gnd VDD3V3 atmpc01_3v3
Xaopac01_3v3_0 LS_3VX2_22|Q AMUX2_3V_0|AOUT analog_out analog_out aopac01_3v3_0|IB  VDD3V3 gnd aopac01_3v3
Xacsoc02_3v3_0 aopac01_3v3_0|IB acsoc02_3v3_0|CS_4U LS_3VX2_19|Q aopac01_3v3_0|IB  acsoc02_3v3_0|CS_8U gnd VDD3V3 acsoc02_3v3
XLS_3VX2_22 LS_3VX2_22|A LS_3VX2_22|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_19 LS_3VX2_19|A LS_3VX2_19|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XBU_3VX2_73 BU_3VX2_73|A BU_3VX2_73|Q gnd vdd BU_3VX2
XAMUX2_3V_0 AMUX4_3V_4|AIN2 AMUX4_3V_4|AIN3 AMUX2_3V_0|AOUT AMUX2_3V_0|SEL vdd VDD3V3 gnd AMUX2_3V__AMUX2_3V 
Xadacc01_3v3_0 AMUX4_3V_4|AIN2 gnd VDD3V3 LS_3VX2_13|Q LS_3VX2_8|Q LS_3VX2_12|Q LS_3VX2_7|Q  LS_3VX2_11|Q LS_3VX2_6|Q LS_3VX2_10|Q LS_3VX2_5|Q LS_3VX2_9|Q LS_3VX2_4|Q LS_3VX2_14|Q  gnd adc_high adc_low VDD3V3 adacc01_3v3
XLS_3VX2_24 LS_3VX2_24|A LS_3VX2_24|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_4 LS_3VX2_4|A LS_3VX2_4|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_5 LS_3VX2_5|A LS_3VX2_5|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_6 LS_3VX2_6|A LS_3VX2_6|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_7 LS_3VX2_7|A LS_3VX2_7|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_8 LS_3VX2_8|A LS_3VX2_8|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_14 LS_3VX2_14|A LS_3VX2_14|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_9 LS_3VX2_9|A LS_3VX2_9|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_10 LS_3VX2_10|A LS_3VX2_10|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_11 LS_3VX2_11|A LS_3VX2_11|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_12 LS_3VX2_12|A LS_3VX2_12|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_13 LS_3VX2_13|A LS_3VX2_13|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
Xraven_soc_0 vdd gnd apllc03_1v8_0|CLK raven_soc_0|ext_clk BU_3VX2_40|Q BU_3VX2_63|Q BU_3VX2_0|Q raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<1> raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<13> raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<15> raven_soc_0|ram_rdata<16> raven_soc_0|ram_rdata<17> raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<31> raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<6> raven_soc_0|gpio_in<7> raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<10> raven_soc_0|gpio_in<11> raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<15> BU_3VX2_43|Q BU_3VX2_44|Q BU_3VX2_45|Q BU_3VX2_46|Q adc0_data<5> BU_3VX2_47|Q BU_3VX2_48|Q BU_3VX2_49|Q BU_3VX2_50|Q BU_3VX2_51|Q BU_3VX2_42|Q BU_3VX2_61|Q BU_3VX2_60|Q BU_3VX2_59|Q BU_3VX2_58|Q BU_3VX2_57|Q BU_3VX2_56|Q BU_3VX2_55|Q BU_3VX2_54|Q BU_3VX2_53|Q BU_3VX2_52|Q BU_3VX2_62|Q BU_3VX2_73|Q BU_3VX2_1|Q BU_3VX2_72|Q BU_3VX2_32|Q BU_3VX2_33|Q BU_3VX2_36|Q BU_3VX2_64|Q BU_3VX2_65|Q BU_3VX2_66|Q BU_3VX2_67|Q BU_3VX2_68|Q BU_3VX2_69|Q BU_3VX2_70|Q BU_3VX2_31|Q BU_3VX2_30|Q BU_3VX2_29|Q BU_3VX2_28|Q BU_3VX2_27|Q BU_3VX2_26|Q BU_3VX2_25|Q BU_3VX2_24|Q BU_3VX2_23|Q BU_3VX2_22|Q BU_3VX2_21|Q BU_3VX2_20|Q BU_3VX2_19|Q BU_3VX2_18|Q BU_3VX2_17|Q BU_3VX2_16|Q BU_3VX2_15|Q BU_3VX2_14|Q BU_3VX2_13|Q BU_3VX2_12|Q BU_3VX2_11|Q BU_3VX2_10|Q BU_3VX2_9|Q BU_3VX2_8|Q BU_3VX2_7|Q BU_3VX2_6|Q BU_3VX2_5|Q BU_3VX2_4|Q BU_3VX2_3|Q BU_3VX2_2|Q BU_3VX2_37|Q BU_3VX2_38|Q BU_3VX2_35|Q raven_soc_0|ser_rx raven_soc_0|irq_pin BU_3VX2_71|Q raven_soc_0|flash_io0_di raven_soc_0|flash_io1_di raven_soc_0|flash_io2_di raven_soc_0|flash_io3_di raven_soc_0|ram_wenb raven_soc_0|ram_addr<0> raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<2> raven_soc_0|ram_addr<3> raven_soc_0|ram_addr<4> raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<22> raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<27> raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<29> raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<31> raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<8> raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<10> raven_soc_0|gpio_out<11> raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<14> raven_soc_0|gpio_out<15> raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<3> raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_outenb<15> LS_3VX2_27|A LS_3VX2_21|A LS_3VX2_20|A AMUX4_3V_0|SEL[0] AMUX4_3V_0|SEL[1] LS_3VX2_17|A LS_3VX2_16|A LS_3VX2_15|A AMUX4_3V_1|SEL[0] AMUX4_3V_1|SEL[1] LS_3VX2_14|A LS_3VX2_4|A LS_3VX2_9|A LS_3VX2_5|A LS_3VX2_10|A LS_3VX2_6|A LS_3VX2_11|A LS_3VX2_7|A LS_3VX2_12|A LS_3VX2_8|A LS_3VX2_13|A AMUX2_3V_0|SEL LS_3VX2_22|A LS_3VX2_19|A LS_3VX2_18|A LS_3VX2_23|A AMUX4_3V_4|SEL[0] AMUX4_3V_4|SEL[1] AMUX4_3V_3|SEL[0] AMUX4_3V_3|SEL[1] LS_3VX2_2|A LS_3VX2_24|A raven_soc_0|ser_tx LS_3VX2_3|A raven_soc_0|flash_csb raven_soc_0|flash_clk raven_soc_0|flash_io0_oeb raven_soc_0|flash_io1_oeb raven_soc_0|flash_io2_oeb raven_soc_0|flash_io3_oeb raven_soc_0|flash_io0_do raven_soc_0|flash_io1_do raven_soc_0|flash_io2_do raven_soc_0|flash_io3_do raven_soc__raven_soc 
Xaadcc01_3v3_0 VDD3V3 BU_3VX2_62|A LS_3VX2_17|Q LS_3VX2_16|Q LS_3VX2_15|Q BU_3VX2_61|A  BU_3VX2_60|A BU_3VX2_59|A BU_3VX2_58|A BU_3VX2_57|A BU_3VX2_56|A BU_3VX2_55|A BU_3VX2_54|A  BU_3VX2_53|A BU_3VX2_52|A AMUX4_3V_1|AOUT adc_high adc_low gnd VDD3V3 gnd aadcc01_3v3
XAMUX4_3V_1 AMUX4_3V_1|AIN1 VDD3V3 AMUX4_3V_4|AIN3 comp_inp AMUX4_3V_1|AOUT AMUX4_3V_1|SEL[1] AMUX4_3V_1|SEL[0] vdd VDD3V3 gnd AMUX4_3V__AMUX4_3V 
Xaadcc01_3v3_1 VDD3V3 BU_3VX2_42|A LS_3VX2_27|Q LS_3VX2_21|Q LS_3VX2_20|Q BU_3VX2_43|A  BU_3VX2_44|A BU_3VX2_45|A BU_3VX2_46|A BU_3VX2_41|A BU_3VX2_47|A BU_3VX2_48|A BU_3VX2_49|A  BU_3VX2_50|A BU_3VX2_51|A AMUX4_3V_0|AOUT adc_high adc_low gnd VDD3V3 gnd aadcc01_3v3
XIN_3VX2_1 IN_3VX2_1|A IN_3VX2_1|Q gnd VDD3V3 IN_3VX2
XAMUX4_3V_0 AMUX4_3V_0|AIN1 vdd AMUX4_3V_4|AIN2 gnd AMUX4_3V_0|AOUT AMUX4_3V_0|SEL[1] AMUX4_3V_0|SEL[0] vdd VDD3V3 gnd AMUX4_3V__AMUX4_3V 
XLS_3VX2_17 LS_3VX2_17|A LS_3VX2_17|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_16 LS_3VX2_16|A LS_3VX2_16|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_15 LS_3VX2_15|A LS_3VX2_15|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XBU_3VX2_62 BU_3VX2_62|A BU_3VX2_62|Q gnd vdd BU_3VX2
XBU_3VX2_61 BU_3VX2_61|A BU_3VX2_61|Q gnd vdd BU_3VX2
XBU_3VX2_60 BU_3VX2_60|A BU_3VX2_60|Q gnd vdd BU_3VX2
XBU_3VX2_59 BU_3VX2_59|A BU_3VX2_59|Q gnd vdd BU_3VX2
XBU_3VX2_58 BU_3VX2_58|A BU_3VX2_58|Q gnd vdd BU_3VX2
XBU_3VX2_57 BU_3VX2_57|A BU_3VX2_57|Q gnd vdd BU_3VX2
XBU_3VX2_56 BU_3VX2_56|A BU_3VX2_56|Q gnd vdd BU_3VX2
XBU_3VX2_55 BU_3VX2_55|A BU_3VX2_55|Q gnd vdd BU_3VX2
XBU_3VX2_54 BU_3VX2_54|A BU_3VX2_54|Q gnd vdd BU_3VX2
XBU_3VX2_53 BU_3VX2_53|A BU_3VX2_53|Q gnd vdd BU_3VX2
XBU_3VX2_52 BU_3VX2_52|A BU_3VX2_52|Q gnd vdd BU_3VX2
XLS_3VX2_27 LS_3VX2_27|A LS_3VX2_27|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_21 LS_3VX2_21|A LS_3VX2_21|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XLS_3VX2_20 LS_3VX2_20|A LS_3VX2_20|Q vdd VDD3V3 gnd LS_3VX2__LS_3VX2 
XBU_3VX2_42 BU_3VX2_42|A BU_3VX2_42|Q gnd vdd BU_3VX2
XBU_3VX2_43 BU_3VX2_43|A BU_3VX2_43|Q gnd vdd BU_3VX2
XBU_3VX2_44 BU_3VX2_44|A BU_3VX2_44|Q gnd vdd BU_3VX2
XBU_3VX2_45 BU_3VX2_45|A BU_3VX2_45|Q gnd vdd BU_3VX2
XBU_3VX2_46 BU_3VX2_46|A BU_3VX2_46|Q gnd vdd BU_3VX2
XBU_3VX2_41 BU_3VX2_41|A adc0_data<5> gnd vdd BU_3VX2
XBU_3VX2_47 BU_3VX2_47|A BU_3VX2_47|Q gnd vdd BU_3VX2
XBU_3VX2_48 BU_3VX2_48|A BU_3VX2_48|Q gnd vdd BU_3VX2
XBU_3VX2_49 BU_3VX2_49|A BU_3VX2_49|Q gnd vdd BU_3VX2
XBU_3VX2_50 BU_3VX2_50|A BU_3VX2_50|Q gnd vdd BU_3VX2
XBU_3VX2_51 BU_3VX2_51|A BU_3VX2_51|Q gnd vdd BU_3VX2
Xapllc03_1v8_0 BU_3VX2_72|Q apllc03_1v8_0|B_VCO apllc03_1v8_0|B_CP vdd gnd BU_3VX2_23|Q  BU_3VX2_24|Q BU_3VX2_25|Q BU_3VX2_26|Q apllc03_1v8_0|VCO_IN apllc03_1v8_0|CLK gnd  vdd BU_3VX2_29|Q BU_3VX2_28|Q apllc03_1v8
Xacsoc04_1v8_0 apllc03_1v8_0|B_CP BU_3VX2_27|Q vdd gnd apllc03_1v8_0|B_VCO apllc03_1v8_0|B_VCO  apllc03_1v8_0|B_CP acsoc04_1v8
XBU_3VX2_72 BU_3VX2_72|A BU_3VX2_72|Q gnd vdd BU_3VX2
C0 AMUX4_3V_1|SEL[1] BU_3VX2_52|Q 63.88fF
C1 AMUX4_3V_3|SEL[1] apllc03_1v8_0|CLK 33.38fF
C2 BU_3VX2_22|A raven_soc_0|flash_csb 2.12fF
C3 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<6> 0.86fF
C4 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<1> 3.58fF
C5 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<11> 22.21fF
C6 BU_3VX2_9|A BU_3VX2_9|Q 0.08fF
C7 LS_3VX2_7|A LS_3VX2_19|A 0.01fF
C8 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<3> 3.52fF
C9 BU_3VX2_31|A raven_soc_0|gpio_in<13> 0.01fF
C10 BU_3VX2_0|Q raven_soc_0|ram_rdata<27> 0.02fF
C11 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<9> 0.28fF
C12 BU_3VX2_13|A VDD3V3 0.53fF
C13 VDD raven_padframe_0|FILLER20F_6|GNDR 0.16fF
C14 LS_3VX2_7|A BU_3VX2_52|Q 9.34fF
C15 adc_high comp_inp 2.71fF
C16 raven_soc_0|ram_wdata<24> raven_soc_0|ram_addr<0> 0.08fF
C17 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<17> 5.90fF
C18 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<16> 5.13fF
C19 LS_3VX2_18|A AMUX4_3V_4|SEL[0] 1.23fF
C20 BU_3VX2_61|Q BU_3VX2_60|Q 233.85fF
C21 LS_3VX2_15|A BU_3VX2_58|Q 25.91fF
C22 BU_3VX2_62|Q BU_3VX2_59|Q 38.82fF
C23 BU_3VX2_46|A BU_3VX2_45|Q 0.15fF
C24 BU_3VX2_46|Q adc0_data<5> 222.29fF
C25 raven_padframe_0|FILLER10F_0|GNDR raven_padframe_0|FILLER10F_0|VDDO 0.09fF
C26 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<12> 0.19fF
C27 raven_soc_0|gpio_in<1> BU_3VX2_23|Q 0.01fF
C28 LS_3VX2_2|Q LS_3VX2_2|A 0.05fF
C29 BU_3VX2_19|A raven_soc_0|flash_io0_di 0.01fF
C30 BU_3VX2_1|A BU_3VX2_32|Q 0.03fF
C31 BU_3VX2_17|A raven_soc_0|flash_io3_do 0.01fF
C32 BU_3VX2_4|A raven_soc_0|flash_io0_do 0.01fF
C33 BU_3VX2_16|A raven_soc_0|flash_io3_oeb 0.01fF
C34 raven_padframe_0|ICFC_1|VDD3 raven_padframe_0|ICFC_1|GNDR 0.16fF
C35 raven_padframe_0|BT4FC_0|VDD3 raven_padframe_0|BT4FC_0|GNDO 0.07fF
C36 raven_padframe_0|FILLER40F_0|VDDR raven_padframe_0|FILLER40F_0|GNDO 0.13fF
C37 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<7> 2.40fF
C38 BU_3VX2_29|A raven_soc_0|flash_io3_oeb 5.88fF
C39 adc_low AMUX4_3V_1|SEL[1] 0.05fF
C40 LS_3VX2_5|A BU_3VX2_59|Q 9.13fF
C41 IN_3VX2_1|A BU_3VX2_28|Q 202.58fF
C42 raven_soc_0|gpio_outenb<10> BU_3VX2_26|Q 0.01fF
C43 raven_soc_0|gpio_pullup<9> BU_3VX2_27|Q 0.01fF
C44 raven_soc_0|gpio_pullup<12> BU_3VX2_29|Q 0.01fF
C45 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<4> 1.07fF
C46 BU_3VX2_68|A BU_3VX2_0|A 0.44fF
C47 BU_3VX2_10|A IN_3VX2_1|A 0.01fF
C48 BU_3VX2_2|A BU_3VX2_29|A 0.01fF
C49 IN_3VX2_1|A raven_soc_0|gpio_pulldown<12> 0.01fF
C50 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<14> 3.34fF
C51 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<5> 0.75fF
C52 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<0> 0.09fF
C53 LS_3VX2_3|A raven_soc_0|gpio_pullup<11> 0.01fF
C54 BU_3VX2_35|A raven_soc_0|flash_io2_di 0.11fF
C55 BU_3VX2_0|Q raven_soc_0|gpio_pulldown<4> 0.01fF
C56 BU_3VX2_25|A raven_soc_0|flash_io1_di 0.01fF
C57 BU_3VX2_37|A raven_soc_0|flash_io3_oeb 0.01fF
C58 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<3> 0.01fF
C59 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<5> 0.01fF
C60 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<15> 33.09fF
C61 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<11> 7.93fF
C62 raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<6> 9.83fF
C63 raven_soc_0|gpio_out<15> VDD3V3 3.58fF
C64 BU_3VX2_58|A LS_3VX2_17|Q 0.19fF
C65 BU_3VX2_57|A BU_3VX2_62|A 0.21fF
C66 BU_3VX2_59|A LS_3VX2_16|Q 0.32fF
C67 BU_3VX2_60|A LS_3VX2_15|Q 0.81fF
C68 AMUX4_3V_0|SEL[1] BU_3VX2_49|Q 11.21fF
C69 BU_3VX2_49|Q BU_3VX2_51|Q 75.42fF
C70 BU_3VX2_42|A vdd 0.06fF
C71 BU_3VX2_22|A BU_3VX2_20|A 13.09fF
C72 BU_3VX2_2|A BU_3VX2_37|A 29.56fF
C73 raven_padframe_0|FILLER20FC_0|GNDR raven_padframe_0|FILLER20FC_0|GNDO 0.81fF
C74 LOGIC1_3V_2|Q LOGIC0_3V_4|Q 0.31fF
C75 raven_padframe_0|APR00DF_5|GNDR raven_padframe_0|APR00DF_5|VDDO 0.09fF
C76 BU_3VX2_0|A IN_3VX2_1|A 0.57fF
C77 BU_3VX2_3|A BU_3VX2_27|A 0.01fF
C78 raven_padframe_0|BBCUD4F_13|VDDO raven_padframe_0|BBCUD4F_13|GNDO 2.28fF
C79 BU_3VX2_15|A BU_3VX2_27|A 1.70fF
C80 raven_padframe_0|FILLER20F_4|VDDR raven_padframe_0|FILLER20F_4|GNDR 0.68fF
C81 raven_padframe_0|aregc01_3v3_0|m4_0_30133# raven_padframe_0|aregc01_3v3_0|m4_0_29057# 0.01fF
C82 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<4> 0.46fF
C83 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<14> 0.18fF
C84 raven_spi_0|sdo_enb raven_soc_0|gpio_outenb<15> 1.35fF
C85 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<2> 4.68fF
C86 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<4> 0.30fF
C87 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<8> 0.01fF
C88 markings_0|efabless_logo_0|m1_8400_n7350# markings_0|efabless_logo_0|m1_7500_n8250# 0.27fF
C89 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<10> 0.02fF
C90 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<11> 0.01fF
C91 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<8> 5.60fF
C92 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<20> 0.16fF
C93 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<13> 0.73fF
C94 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<6> 0.01fF
C95 raven_soc_0|gpio_outenb<13> raven_soc_0|ext_clk 0.01fF
C96 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<9> 92.13fF
C97 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<15> 0.02fF
C98 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<0> 0.01fF
C99 LS_3VX2_23|A VDD3V3 0.52fF
C100 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<1> 0.02fF
C101 LS_3VX2_22|A LS_3VX2_15|A 0.02fF
C102 raven_soc_0|gpio_in<5> VDD3V3 0.07fF
C103 LS_3VX2_18|A vdd 1.77fF
C104 BU_3VX2_17|Q BU_3VX2_27|Q 3.52fF
C105 BU_3VX2_21|A raven_soc_0|flash_csb 1.89fF
C106 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<7> 0.68fF
C107 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<15> 1.41fF
C108 BU_3VX2_12|A raven_soc_0|flash_io3_do 0.01fF
C109 VDD raven_padframe_0|VDDORPADF_2|GNDO 0.07fF
C110 raven_soc_0|gpio_pullup<0> vdd 0.22fF
C111 VDD raven_padframe_0|BBCUD4F_7|GNDR 0.16fF
C112 BU_3VX2_0|Q BU_3VX2_7|Q 0.01fF
C113 BU_3VX2_0|Q BU_3VX2_6|Q 0.01fF
C114 adc_high vdd 0.15fF
C115 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_out<14> 0.02fF
C116 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<20> 4.40fF
C117 raven_soc_0|ram_rdata<21> raven_soc_0|ram_addr<3> 1.02fF
C118 raven_soc_0|ram_rdata<7> raven_soc_0|ram_addr<2> 0.04fF
C119 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<30> 6.29fF
C120 raven_soc_0|ram_rdata<5> raven_soc_0|ram_addr<4> 0.24fF
C121 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<8> 6.02fF
C122 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<9> 2.60fF
C123 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_out<10> 0.01fF
C124 BU_3VX2_14|Q BU_3VX2_3|Q 3.07fF
C125 AMUX4_3V_1|SEL[1] BU_3VX2_58|Q 12.22fF
C126 raven_soc_0|ram_rdata<19> apllc03_1v8_0|CLK 0.01fF
C127 raven_padframe_0|ICFC_2|GNDR raven_padframe_0|ICFC_2|GNDO 0.81fF
C128 raven_padframe_0|axtoc02_3v3_0|m4_55000_0# raven_padframe_0|axtoc02_3v3_0|GNDO 2.48fF
C129 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<12> 0.17fF
C130 BU_3VX2_23|A vdd 0.06fF
C131 LS_3VX2_9|A AMUX4_3V_1|SEL[0] 33.40fF
C132 BU_3VX2_67|A BU_3VX2_64|Q 0.02fF
C133 LS_3VX2_3|Q raven_soc_0|flash_io3_oeb 0.01fF
C134 LS_3VX2_7|A BU_3VX2_58|Q 0.01fF
C135 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<8> 0.51fF
C136 IN_3VX2_1|A BU_3VX2_44|Q 11.03fF
C137 IN_3VX2_1|A comp_inp 2.28fF
C138 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<7> 15.18fF
C139 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<14> 17.57fF
C140 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<15> 313.44fF
C141 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<8> 17.68fF
C142 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<13> 0.51fF
C143 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<6> 0.19fF
C144 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<12> 59.72fF
C145 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<10> 19.33fF
C146 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<15> 0.02fF
C147 BU_3VX2_0|Q raven_soc_0|flash_io2_di 0.01fF
C148 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pullup<5> 0.02fF
C149 BU_3VX2_2|A LS_3VX2_3|Q 0.01fF
C150 LS_3VX2_7|Q LS_3VX2_4|Q 0.61fF
C151 BU_3VX2_31|A raven_soc_0|gpio_outenb<1> 0.01fF
C152 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_in<2> 7.11fF
C153 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<6> 0.01fF
C154 LOGIC0_3V_4|Q raven_soc_0|flash_io3_oeb 0.01fF
C155 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<10> 0.48fF
C156 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<13> 1.94fF
C157 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pullup<6> 0.02fF
C158 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pullup<14> 48.26fF
C159 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pullup<13> 0.01fF
C160 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<5> 0.13fF
C161 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<13> 0.01fF
C162 raven_soc_0|gpio_pullup<15> BU_3VX2_71|Q 0.01fF
C163 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<13> 0.19fF
C164 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<1> 0.01fF
C165 AMUX2_3V_0|SEL BU_3VX2_62|Q 0.01fF
C166 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<26> 0.19fF
C167 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<3> 0.02fF
C168 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<2> 1.29fF
C169 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<12> 0.01fF
C170 BU_3VX2_16|Q BU_3VX2_6|Q 6.59fF
C171 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<15> 4.17fF
C172 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<25> 0.39fF
C173 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<17> 8.57fF
C174 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<14> 15.77fF
C175 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<13> 20.81fF
C176 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<2> 0.09fF
C177 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<8> 0.01fF
C178 BU_3VX2_68|Q BU_3VX2_8|Q 3.81fF
C179 BU_3VX2_16|Q BU_3VX2_7|Q 3.83fF
C180 BU_3VX2_21|Q BU_3VX2_68|Q 25.25fF
C181 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<14> 7.63fF
C182 BU_3VX2_65|Q BU_3VX2_22|Q 4.52fF
C183 BU_3VX2_64|Q BU_3VX2_10|Q 0.03fF
C184 raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<13> 2.13fF
C185 BU_3VX2_12|Q BU_3VX2_69|Q 0.53fF
C186 BU_3VX2_30|Q BU_3VX2_7|Q 6.38fF
C187 BU_3VX2_2|Q BU_3VX2_64|Q 0.67fF
C188 BU_3VX2_13|Q BU_3VX2_5|Q 7.18fF
C189 BU_3VX2_31|Q BU_3VX2_67|Q 0.66fF
C190 BU_3VX2_43|Q BU_3VX2_48|Q 20.85fF
C191 BU_3VX2_21|A BU_3VX2_20|A 36.61fF
C192 raven_padframe_0|CORNERESDF_3|VDDO raven_padframe_0|CORNERESDF_3|GNDO 2.28fF
C193 BU_3VX2_10|A BU_3VX2_25|A 0.01fF
C194 BU_3VX2_8|A BU_3VX2_17|A 1.32fF
C195 BU_3VX2_19|A BU_3VX2_5|A 0.01fF
C196 raven_padframe_0|FILLER20F_6|VDDR raven_padframe_0|FILLER20F_6|GNDO 0.13fF
C197 raven_padframe_0|FILLER20F_6|GNDR raven_padframe_0|FILLER20F_6|VDDO 0.09fF
C198 BU_3VX2_65|A BU_3VX2_36|A 8.33fF
C199 LS_3VX2_5|A AMUX2_3V_0|SEL 10.14fF
C200 raven_soc_0|gpio_pulldown<11> BU_3VX2_0|Q 0.01fF
C201 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<5> 0.13fF
C202 raven_soc_0|gpio_pulldown<8> LS_3VX2_3|A 0.01fF
C203 LS_3VX2_22|A AMUX4_3V_1|SEL[1] 6.86fF
C204 raven_soc_0|ram_wdata<31> vdd 1.06fF
C205 BU_3VX2_25|A BU_3VX2_0|A 0.01fF
C206 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<4> 0.01fF
C207 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<11> 0.84fF
C208 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<11> 0.01fF
C209 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<13> 10.52fF
C210 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<9> 1.08fF
C211 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<5> 0.03fF
C212 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<11> 14.37fF
C213 markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# markings_0|product_name_0|_alphabet_V_0|m2_0_560# 0.11fF
C214 BU_3VX2_2|A BU_3VX2_38|Q 0.03fF
C215 BU_3VX2_68|A vdd 0.22fF
C216 LS_3VX2_7|A LS_3VX2_22|A 14.75fF
C217 BU_3VX2_4|A BU_3VX2_5|Q 0.03fF
C218 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<17> 0.05fF
C219 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<29> 30.18fF
C220 raven_soc_0|flash_io3_di raven_soc_0|flash_io2_di 393.00fF
C221 raven_soc_0|flash_io0_oeb raven_soc_0|flash_io0_do 66.44fF
C222 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<1> 0.05fF
C223 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<16> 30.75fF
C224 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io1_oeb 120.50fF
C225 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<31> 4.28fF
C226 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<22> 0.12fF
C227 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<13> 0.23fF
C228 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<15> 1.95fF
C229 raven_soc_0|ram_rdata<8> raven_soc_0|ram_addr<0> 0.05fF
C230 BU_3VX2_1|Q BU_3VX2_32|Q 0.27fF
C231 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<24> 0.01fF
C232 BU_3VX2_62|Q BU_3VX2_61|Q 123.30fF
C233 LS_3VX2_15|A BU_3VX2_60|Q 59.63fF
C234 raven_padframe_0|GNDORPADF_0|VDDR raven_padframe_0|GNDORPADF_0|VDDO 0.06fF
C235 raven_padframe_0|FILLER20F_2|VDDO raven_padframe_0|FILLER20F_2|GNDO 2.28fF
C236 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<12> 0.53fF
C237 BU_3VX2_2|A raven_soc_0|flash_io1_oeb 0.01fF
C238 BU_3VX2_35|A BU_3VX2_35|Q 0.08fF
C239 LS_3VX2_9|A LS_3VX2_17|A 0.43fF
C240 BU_3VX2_4|A raven_soc_0|flash_io1_di 0.07fF
C241 IN_3VX2_1|Q BU_3VX2_52|Q 0.01fF
C242 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<9> 0.01fF
C243 raven_padframe_0|FILLER20FC_0|VDD3 raven_padframe_0|FILLER20FC_0|GNDO 0.07fF
C244 raven_padframe_0|VDDPADFC_0|VDDR raven_padframe_0|VDDPADFC_0|GNDO 0.13fF
C245 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<7> 0.25fF
C246 LS_3VX2_8|A BU_3VX2_54|Q 6.23fF
C247 raven_soc_0|gpio_in<4> BU_3VX2_40|Q 0.01fF
C248 IN_3VX2_1|A vdd 1.95fF
C249 BU_3VX2_14|A BU_3VX2_15|Q 0.03fF
C250 LS_3VX2_5|A BU_3VX2_61|Q 0.01fF
C251 LS_3VX2_13|A BU_3VX2_73|Q 17.66fF
C252 raven_soc_0|gpio_pullup<10> BU_3VX2_26|Q 0.01fF
C253 raven_soc_0|gpio_pullup<9> BU_3VX2_25|Q 0.01fF
C254 raven_soc_0|gpio_pulldown<9> BU_3VX2_27|Q 0.01fF
C255 raven_soc_0|gpio_outenb<0> BU_3VX2_29|Q 0.01fF
C256 BU_3VX2_8|A BU_3VX2_12|A 3.17fF
C257 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<7> 0.01fF
C258 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<5> 1.34fF
C259 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<3> 0.01fF
C260 BU_3VX2_72|A BU_3VX2_72|Q 0.09fF
C261 raven_soc_0|ext_clk raven_soc_0|gpio_in<8> 0.01fF
C262 BU_3VX2_40|Q raven_soc_0|gpio_in<7> 0.01fF
C263 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<12> 0.02fF
C264 raven_soc_0|gpio_in<6> VDD3V3 0.07fF
C265 BU_3VX2_53|A BU_3VX2_59|A 0.59fF
C266 BU_3VX2_52|A BU_3VX2_60|A 0.36fF
C267 BU_3VX2_54|A BU_3VX2_58|A 1.07fF
C268 BU_3VX2_55|A BU_3VX2_57|A 3.29fF
C269 VDD3V3 LS_3VX2_15|Q 0.35fF
C270 raven_soc_0|irq_pin BU_3VX2_55|Q 0.01fF
C271 raven_soc_0|gpio_in<1> BU_3VX2_31|A 0.01fF
C272 BU_3VX2_48|Q BU_3VX2_50|Q 75.11fF
C273 BU_3VX2_38|A BU_3VX2_35|A 30.16fF
C274 BU_3VX2_71|A BU_3VX2_18|A 0.01fF
C275 IN_3VX2_1|Q adc_low 0.05fF
C276 BU_3VX2_40|A IN_3VX2_1|A 0.12fF
C277 IN_3VX2_1|A raven_soc_0|gpio_in<2> 0.01fF
C278 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<15> 0.46fF
C279 markings_0|efabless_logo_0|m1_8400_n4650# markings_0|efabless_logo_0|m1_8700_n6150# 0.23fF
C280 raven_soc_0|gpio_out<3> BU_3VX2_71|Q 0.01fF
C281 raven_soc_0|gpio_out<10> VDD3V3 0.07fF
C282 raven_soc_0|flash_io2_di raven_soc_0|irq_pin 0.01fF
C283 raven_soc_0|gpio_pullup<13> raven_soc_0|ext_clk 0.01fF
C284 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<13> 0.02fF
C285 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<14> 0.02fF
C286 BU_3VX2_21|Q BU_3VX2_24|Q 21.37fF
C287 BU_3VX2_8|Q BU_3VX2_24|Q 2.04fF
C288 BU_3VX2_20|Q BU_3VX2_23|Q 13.17fF
C289 BU_3VX2_12|Q BU_3VX2_29|Q 0.84fF
C290 BU_3VX2_13|Q BU_3VX2_28|Q 0.54fF
C291 BU_3VX2_66|Q BU_3VX2_23|Q 0.41fF
C292 BU_3VX2_17|Q BU_3VX2_25|Q 4.39fF
C293 BU_3VX2_38|Q apllc03_1v8_0|CLK 0.01fF
C294 BU_3VX2_67|Q apllc03_1v8_0|CLK 0.93fF
C295 BU_3VX2_0|A aporc02_3v3_0|PORB 0.65fF
C296 BU_3VX2_67|A BU_3VX2_33|A 1.39fF
C297 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<7> 0.01fF
C298 LS_3VX2_5|Q VDD3V3 0.16fF
C299 BU_3VX2_70|A BU_3VX2_67|Q 0.02fF
C300 BU_3VX2_26|A raven_soc_0|ext_clk 0.01fF
C301 LS_3VX2_24|A BU_3VX2_50|Q 7.88fF
C302 BU_3VX2_0|Q BU_3VX2_35|Q 0.01fF
C303 raven_soc_0|ser_rx BU_3VX2_73|Q 0.01fF
C304 LS_3VX2_4|A BU_3VX2_54|Q 20.43fF
C305 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<18> 8.02fF
C306 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<14> 6.58fF
C307 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<21> 0.01fF
C308 raven_soc_0|ram_addr<0> raven_soc_0|ram_rdata<16> 0.39fF
C309 raven_soc_0|flash_io0_di BU_3VX2_27|Q 0.01fF
C310 raven_soc_0|flash_io0_do BU_3VX2_29|Q 0.01fF
C311 AMUX4_3V_1|SEL[1] BU_3VX2_60|Q 9.63fF
C312 raven_soc_0|flash_io1_oeb apllc03_1v8_0|CLK 0.01fF
C313 raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# raven_padframe_0|axtoc02_3v3_0|VDDO 0.07fF
C314 markings_0|manufacturer_0|_alphabet_S_0|m2_32_224# markings_0|manufacturer_0|_alphabet_E_2|m2_0_0# 0.14fF
C315 abgpc01_3v3_0|VBGVTN VDD3V3 0.05fF
C316 LS_3VX2_10|A raven_soc_0|ser_tx 0.01fF
C317 BU_3VX2_63|A raven_soc_0|flash_io2_di 0.01fF
C318 LS_3VX2_7|A BU_3VX2_60|Q 0.01fF
C319 BU_3VX2_11|A raven_soc_0|ext_clk 0.01fF
C320 IN_3VX2_1|A raven_soc_0|gpio_in<11> 0.01fF
C321 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<12> 166.14fF
C322 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<9> 0.91fF
C323 LS_3VX2_6|A BU_3VX2_55|Q 8.52fF
C324 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<8> 5.26fF
C325 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<14> 34.71fF
C326 raven_soc_0|gpio_out<7> BU_3VX2_40|Q 0.01fF
C327 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<10> 10.48fF
C328 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<7> 42.94fF
C329 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<13> 7.49fF
C330 raven_soc_0|gpio_out<9> VDD3V3 0.07fF
C331 raven_soc_0|gpio_in<3> VDD3V3 0.44fF
C332 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<6> 18.34fF
C333 raven_soc_0|gpio_out<5> raven_soc_0|ext_clk 0.01fF
C334 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<15> 0.02fF
C335 raven_padframe_0|BBCUD4F_3|VDDR raven_padframe_0|BBCUD4F_3|GNDR 0.68fF
C336 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<0> 0.01fF
C337 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<19> 0.02fF
C338 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<20> 12.21fF
C339 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<23> 0.04fF
C340 BU_3VX2_10|A BU_3VX2_4|A 1.98fF
C341 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<8> 0.01fF
C342 LS_3VX2_10|A LS_3VX2_24|A 8.72fF
C343 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<7> 0.01fF
C344 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<2> 7.61fF
C345 BU_3VX2_3|A BU_3VX2_37|Q 0.03fF
C346 IN_3VX2_1|Q BU_3VX2_58|Q 0.01fF
C347 LS_3VX2_11|A BU_3VX2_59|Q 0.04fF
C348 BU_3VX2_25|A vdd 0.06fF
C349 IN_3VX2_1|A raven_soc_0|gpio_outenb<9> 0.01fF
C350 raven_soc_0|ram_wenb raven_soc_0|ram_addr<7> 0.01fF
C351 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pullup<13> 0.16fF
C352 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<13> 7.43fF
C353 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<8> 0.21fF
C354 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<10> 0.15fF
C355 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pullup<14> 35.77fF
C356 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pulldown<7> 0.02fF
C357 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pullup<6> 0.02fF
C358 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<5> 0.01fF
C359 BU_3VX2_33|A raven_soc_0|flash_clk 0.01fF
C360 raven_soc_0|gpio_pulldown<14> BU_3VX2_29|Q 0.01fF
C361 BU_3VX2_63|Q BU_3VX2_27|Q 2.30fF
C362 raven_soc_0|gpio_pulldown<15> BU_3VX2_23|Q 0.01fF
C363 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<16> 16.82fF
C364 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<18> 6.70fF
C365 BU_3VX2_19|Q BU_3VX2_68|Q 0.01fF
C366 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<8> 16.57fF
C367 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<2> 2.36fF
C368 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<25> 3.15fF
C369 BU_3VX2_68|Q BU_3VX2_18|Q 5.45fF
C370 BU_3VX2_5|Q BU_3VX2_69|Q 7.94fF
C371 AMUX4_3V_3|SEL[0] BU_3VX2_7|Q 0.03fF
C372 BU_3VX2_31|Q BU_3VX2_65|Q 0.50fF
C373 BU_3VX2_64|Q BU_3VX2_33|Q 0.51fF
C374 LS_3VX2_21|Q BU_3VX2_42|Q 1.07fF
C375 VDD raven_padframe_0|BT4F_2|VDDR 0.71fF
C376 raven_padframe_0|FILLER20F_1|GNDR raven_padframe_0|FILLER20F_1|VDDO 0.09fF
C377 BU_3VX2_0|A BU_3VX2_4|A 0.09fF
C378 LS_3VX2_14|A LS_3VX2_8|A 53.27fF
C379 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<0> 6.19fF
C380 BU_3VX2_19|A BU_3VX2_13|A 2.98fF
C381 raven_padframe_0|BBCUD4F_7|GNDR raven_padframe_0|BBCUD4F_7|VDDO 0.09fF
C382 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<15> 0.01fF
C383 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<13> 0.01fF
C384 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<8> 0.01fF
C385 raven_soc_0|ram_addr<5> vdd 0.51fF
C386 raven_soc_0|ram_wdata<19> vdd 1.03fF
C387 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<6> 0.49fF
C388 raven_padframe_0|BT4F_2|VDDR LOGIC0_3V_4|Q 0.01fF
C389 aopac01_3v3_0|IB AMUX2_3V_0|AOUT 0.44fF
C390 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<3> 43.30fF
C391 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<1> 0.52fF
C392 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<6> 0.01fF
C393 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<11> 0.01fF
C394 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<7> 49.46fF
C395 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<5> 0.02fF
C396 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<9> 0.18fF
C397 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<6> 0.14fF
C398 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<11> 9.33fF
C399 raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<3> 10.30fF
C400 raven_soc_0|flash_io1_di raven_soc_0|flash_io0_oeb 19.86fF
C401 BU_3VX2_66|Q BU_3VX2_4|Q 2.57fF
C402 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<13> 4.17fF
C403 raven_soc_0|flash_io2_do raven_soc_0|flash_io0_do 131.09fF
C404 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<4> 21.95fF
C405 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<1> 0.34fF
C406 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<27> 25.25fF
C407 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<10> 0.15fF
C408 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<17> 0.04fF
C409 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<24> 0.15fF
C410 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<19> 0.32fF
C411 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io0_di 16.34fF
C412 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<2> 12.95fF
C413 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<31> 0.02fF
C414 raven_soc_0|ram_rdata<22> raven_soc_0|ram_addr<0> 5.19fF
C415 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<25> 18.37fF
C416 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<22> 0.01fF
C417 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<29> 3.08fF
C418 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<21> 0.01fF
C419 raven_soc_0|flash_io3_do raven_soc_0|flash_clk 16.56fF
C420 BU_3VX2_36|Q BU_3VX2_22|Q 0.38fF
C421 raven_soc_0|flash_clk AMUX4_3V_4|AIN3 9.29fF
C422 LS_3VX2_15|A BU_3VX2_62|Q 169.60fF
C423 raven_padframe_0|FILLER20F_5|GNDR raven_padframe_0|FILLER20F_5|VDDO 0.09fF
C424 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<0> 27.40fF
C425 raven_spi_0|SDO raven_soc_0|flash_io2_di 1.05fF
C426 BU_3VX2_6|A raven_soc_0|flash_io0_di 0.03fF
C427 BU_3VX2_9|A raven_soc_0|flash_io3_do 0.01fF
C428 BU_3VX2_38|A raven_soc_0|flash_io3_di 0.01fF
C429 LS_3VX2_8|A BU_3VX2_56|Q 2.47fF
C430 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<6> 0.01fF
C431 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<3> 4.47fF
C432 LS_3VX2_5|A LS_3VX2_15|A 0.02fF
C433 raven_padframe_0|BBCUD4F_13|VDDR raven_padframe_0|BBCUD4F_13|GNDR 0.68fF
C434 raven_soc_0|gpio_pulldown<13> apllc03_1v8_0|CLK 0.35fF
C435 raven_soc_0|gpio_pullup<3> vdd 0.33fF
C436 BU_3VX2_0|Q BU_3VX2_23|Q 0.02fF
C437 raven_soc_0|gpio_pulldown<10> BU_3VX2_29|Q 0.01fF
C438 raven_soc_0|gpio_pulldown<9> BU_3VX2_25|Q 0.01fF
C439 LS_3VX2_14|A LS_3VX2_4|A 9.57fF
C440 raven_soc_0|gpio_out<4> BU_3VX2_0|Q 0.01fF
C441 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<5> 0.72fF
C442 aopac01_3v3_0|IB LS_3VX2_22|A 0.01fF
C443 AMUX4_3V_4|AOUT comp_inp 0.02fF
C444 BU_3VX2_63|Q raven_soc_0|flash_io2_oeb 0.03fF
C445 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<10> 5.34fF
C446 raven_soc_0|gpio_pulldown<0> BU_3VX2_23|Q 0.01fF
C447 raven_soc_0|gpio_pullup<1> apllc03_1v8_0|CLK 0.01fF
C448 raven_soc_0|gpio_out<2> BU_3VX2_27|Q 0.01fF
C449 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_2|PO 0.04fF
C450 BU_3VX2_24|A BU_3VX2_18|A 3.69fF
C451 raven_soc_0|ext_clk VDD3V3 7.09fF
C452 raven_soc_0|irq_pin BU_3VX2_57|Q 0.01fF
C453 VDD3V3 BU_3VX2_52|A 0.05fF
C454 LS_3VX2_21|Q BU_3VX2_42|A 1.87fF
C455 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<2> 9.01fF
C456 VDD raven_padframe_0|FILLER20F_1|VDDR 0.71fF
C457 raven_padframe_0|POWERCUTVDD3FC_0|GNDR raven_padframe_0|POWERCUTVDD3FC_0|VDDO 0.09fF
C458 raven_padframe_0|BBCUD4F_3|GNDR raven_padframe_0|BBCUD4F_3|GNDO 0.81fF
C459 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<4> 0.87fF
C460 BU_3VX2_31|A raven_soc_0|gpio_pullup<7> 0.01fF
C461 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<11> 0.01fF
C462 raven_soc_0|gpio_outenb<2> LS_3VX2_3|A 0.01fF
C463 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<3> 1.79fF
C464 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<14> 0.01fF
C465 raven_padframe_0|BBCUD4F_14|VDDR raven_padframe_0|BBCUD4F_14|VDDO 0.06fF
C466 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<11> 0.01fF
C467 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pullup<5> 1.77fF
C468 BU_3VX2_16|Q BU_3VX2_23|Q 5.29fF
C469 BU_3VX2_13|Q vdd 1.42fF
C470 BU_3VX2_19|Q BU_3VX2_24|Q 8.31fF
C471 BU_3VX2_73|Q BU_3VX2_72|Q 19.81fF
C472 BU_3VX2_6|Q BU_3VX2_26|Q 0.01fF
C473 AMUX4_3V_4|AIN2 BU_3VX2_53|Q 0.01fF
C474 BU_3VX2_30|Q BU_3VX2_23|Q 6.84fF
C475 BU_3VX2_18|Q BU_3VX2_24|Q 7.69fF
C476 BU_3VX2_68|Q BU_3VX2_27|Q 3.77fF
C477 BU_3VX2_69|Q BU_3VX2_28|Q 0.50fF
C478 BU_3VX2_7|Q BU_3VX2_26|Q 0.02fF
C479 BU_3VX2_5|Q BU_3VX2_29|Q 0.01fF
C480 BU_3VX2_65|Q apllc03_1v8_0|CLK 0.96fF
C481 BU_3VX2_54|Q vdd 1.62fF
C482 VDD raven_padframe_0|FILLER10F_0|VDDR 0.71fF
C483 raven_padframe_0|FILLER20F_1|VDDR LOGIC0_3V_4|Q 0.01fF
C484 raven_padframe_0|ICFC_1|VDDR LOGIC0_3V_4|Q 0.01fF
C485 raven_soc_0|gpio_pullup<2> IN_3VX2_1|A 0.01fF
C486 LS_3VX2_11|A AMUX2_3V_0|SEL 14.89fF
C487 LOGIC0_3V_4|Q raven_spi_0|sdo_enb 0.75fF
C488 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<9> 0.01fF
C489 LS_3VX2_24|A BU_3VX2_48|Q 6.25fF
C490 LS_3VX2_4|A BU_3VX2_56|Q 13.17fF
C491 raven_soc_0|gpio_pulldown<3> raven_soc_0|gpio_pulldown<6> 1.22fF
C492 raven_soc_0|ram_wdata<29> raven_soc_0|ram_rdata<16> 0.02fF
C493 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<16> 0.01fF
C494 LS_3VX2_2|A LS_3VX2_18|A 4.74fF
C495 AMUX4_3V_1|SEL[1] BU_3VX2_62|Q 9.06fF
C496 BU_3VX2_51|A vdd 0.16fF
C497 raven_soc_0|flash_io3_di BU_3VX2_23|Q 0.01fF
C498 raven_soc_0|flash_io0_di BU_3VX2_25|Q 0.01fF
C499 raven_soc_0|flash_io2_di BU_3VX2_26|Q 0.01fF
C500 raven_soc_0|flash_io0_oeb BU_3VX2_28|Q 13.33fF
C501 raven_soc_0|flash_io1_di BU_3VX2_29|Q 0.01fF
C502 BU_3VX2_59|A BU_3VX2_58|Q 0.03fF
C503 raven_padframe_0|ICF_0|VDDO raven_padframe_0|ICF_0|GNDO 2.28fF
C504 raven_padframe_0|FILLER10F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C505 raven_padframe_0|aregc01_3v3_1|m4_92500_0# raven_padframe_0|aregc01_3v3_1|GNDO 1.24fF
C506 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<8> 0.01fF
C507 markings_0|date_0|_alphabet_0_0|m2_0_208# markings_0|manufacturer_0|_alphabet_E_2|m2_0_0# 0.15fF
C508 VDD raven_soc_0|gpio_in<15> 0.20fF
C509 BU_3VX2_10|A raven_soc_0|flash_io0_oeb 0.01fF
C510 BU_3VX2_4|A vdd 0.51fF
C511 LS_3VX2_24|A raven_soc_0|ser_tx 0.01fF
C512 BU_3VX2_65|A VDD3V3 0.02fF
C513 BU_3VX2_28|A raven_soc_0|flash_io3_do 3.43fF
C514 LS_3VX2_7|A BU_3VX2_62|Q 0.01fF
C515 BU_3VX2_33|A BU_3VX2_33|Q 0.08fF
C516 LS_3VX2_6|A BU_3VX2_57|Q 7.85fF
C517 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<9> 0.02fF
C518 raven_soc_0|gpio_outenb<7> BU_3VX2_40|Q 0.67fF
C519 LS_3VX2_5|A AMUX4_3V_1|SEL[1] 33.29fF
C520 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<7> 2.41fF
C521 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<6> 1.22fF
C522 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<8> 3.59fF
C523 raven_soc_0|gpio_outenb<6> raven_soc_0|ext_clk 0.01fF
C524 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<13> 11.54fF
C525 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<12> 61.79fF
C526 VDD raven_padframe_0|APR00DF_0|GNDO 0.07fF
C527 raven_soc_0|gpio_outenb<10> VDD3V3 0.07fF
C528 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<28> 9.46fF
C529 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<19> 5.00fF
C530 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<23> 6.74fF
C531 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<20> 10.33fF
C532 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<11> 0.30fF
C533 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<0> 1.53fF
C534 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<14> 0.01fF
C535 BU_3VX2_38|A BU_3VX2_63|A 0.01fF
C536 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<6> 0.01fF
C537 LS_3VX2_7|A LS_3VX2_5|A 23.22fF
C538 BU_3VX2_8|A raven_soc_0|flash_clk 0.01fF
C539 BU_3VX2_5|A raven_soc_0|flash_io2_oeb 0.01fF
C540 LS_3VX2_11|A BU_3VX2_61|Q 0.01fF
C541 LS_3VX2_12|A BU_3VX2_51|Q 4.62fF
C542 IN_3VX2_1|Q BU_3VX2_60|Q 0.01fF
C543 BU_3VX2_0|A raven_soc_0|flash_io0_oeb 3.46fF
C544 AMUX4_3V_4|AOUT vdd 0.43fF
C545 LOGIC0_3V_4|Q raven_soc_0|gpio_in<15> 38.78fF
C546 raven_spi_0|sdo_enb raven_soc_0|flash_io1_oeb 0.48fF
C547 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<8> 0.01fF
C548 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<13> 2.54fF
C549 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_outenb<9> 0.46fF
C550 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pulldown<7> 0.02fF
C551 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<10> 8.71fF
C552 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pulldown<6> 0.58fF
C553 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<8> 63.46fF
C554 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<2> 0.01fF
C555 BU_3VX2_0|Q BU_3VX2_4|Q 0.01fF
C556 BU_3VX2_27|A raven_soc_0|flash_io0_di 0.01fF
C557 VDD raven_padframe_0|axtoc02_3v3_0|GNDO 0.11fF
C558 raven_soc_0|gpio_pulldown<11> BU_3VX2_26|Q 0.01fF
C559 BU_3VX2_63|Q BU_3VX2_25|Q 1.93fF
C560 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<12> 2.46fF
C561 raven_soc_0|ram_wdata<0> raven_soc_0|ram_rdata<12> 0.05fF
C562 BU_3VX2_8|A BU_3VX2_9|A 32.91fF
C563 BU_3VX2_23|A BU_3VX2_7|A 0.01fF
C564 BU_3VX2_6|A BU_3VX2_5|A 21.99fF
C565 VDD raven_padframe_0|GNDORPADF_7|VDDR 0.71fF
C566 BU_3VX2_16|A BU_3VX2_18|A 13.47fF
C567 BU_3VX2_4|A BU_3VX2_40|A 1.14fF
C568 raven_padframe_0|VDDPADF_0|VDDO raven_padframe_0|VDDPADF_0|GNDO 2.28fF
C569 BU_3VX2_68|A BU_3VX2_69|A 25.13fF
C570 BU_3VX2_18|A BU_3VX2_29|A 1.94fF
C571 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_outenb<8> 0.19fF
C572 AMUX2_3V_0|SEL LS_3VX2_21|A 11.45fF
C573 raven_soc_0|flash_io3_do BU_3VX2_33|Q 0.01fF
C574 BU_3VX2_73|Q AMUX4_3V_1|SEL[0] 0.01fF
C575 BU_3VX2_24|A BU_3VX2_71|A 0.01fF
C576 raven_soc_0|ram_wdata<30> vdd 0.84fF
C577 raven_soc_0|irq_pin LS_3VX2_16|A 0.01fF
C578 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<11> 0.01fF
C579 BU_3VX2_3|A BU_3VX2_15|A 0.82fF
C580 BU_3VX2_35|A BU_3VX2_31|A 0.01fF
C581 raven_padframe_0|GNDORPADF_7|VDDR LOGIC0_3V_4|Q 0.01fF
C582 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<4> 0.15fF
C583 BU_3VX2_31|A raven_soc_0|gpio_pulldown<15> 0.01fF
C584 IN_3VX2_1|A raven_soc_0|gpio_outenb<14> 0.01fF
C585 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<8> 0.01fF
C586 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<11> 0.37fF
C587 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<10> 0.70fF
C588 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<5> 0.01fF
C589 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<6> 1.58fF
C590 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<7> 0.01fF
C591 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<9> 87.16fF
C592 acsoc01_3v3_0|CS2_200N VDD3V3 0.02fF
C593 LS_3VX2_12|Q VDD3V3 0.21fF
C594 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<3> 6.81fF
C595 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<9> 12.53fF
C596 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<6> 3.63fF
C597 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<8> 2.38fF
C598 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<31> 0.01fF
C599 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<22> 0.01fF
C600 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<23> 0.01fF
C601 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<24> 3.76fF
C602 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<18> 0.01fF
C603 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<13> 7.66fF
C604 BU_3VX2_6|Q BU_3VX2_11|Q 35.96fF
C605 BU_3VX2_13|Q BU_3VX2_70|Q 36.37fF
C606 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<2> 0.07fF
C607 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<26> 35.75fF
C608 BU_3VX2_16|Q BU_3VX2_4|Q 3.17fF
C609 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<29> 0.19fF
C610 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<25> 0.31fF
C611 raven_soc_0|flash_io2_do raven_soc_0|flash_io1_di 58.38fF
C612 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<15> 4.57fF
C613 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<21> 0.02fF
C614 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<14> 0.01fF
C615 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<25> 0.01fF
C616 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<22> 3.60fF
C617 BU_3VX2_4|Q BU_3VX2_30|Q 2.18fF
C618 BU_3VX2_37|Q BU_3VX2_17|Q 3.59fF
C619 BU_3VX2_11|Q BU_3VX2_7|Q 10.06fF
C620 BU_3VX2_36|Q BU_3VX2_31|Q 0.01fF
C621 BU_3VX2_24|Q BU_3VX2_27|Q 72.66fF
C622 BU_3VX2_28|Q BU_3VX2_29|Q 346.91fF
C623 apllc03_1v8_0|B_VCO apllc03_1v8_0|B_CP 26.31fF
C624 apllc03_1v8_0|CLK BU_3VX2_72|Q 0.03fF
C625 raven_padframe_0|BBCUD4F_15|VDDO raven_padframe_0|BBCUD4F_15|GNDO 2.28fF
C626 raven_padframe_0|FILLER50F_1|GNDR raven_padframe_0|FILLER50F_1|GNDO 0.81fF
C627 LOGIC0_3V_4|Q raven_soc_0|gpio_out<13> 0.01fF
C628 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<10> 0.01fF
C629 AMUX4_3V_1|AIN1 comp_inp 1.59fF
C630 LS_3VX2_14|A vdd 2.90fF
C631 raven_soc_0|gpio_pulldown<12> BU_3VX2_29|Q 0.01fF
C632 raven_soc_0|gpio_pulldown<5> vdd 0.44fF
C633 VDD raven_padframe_0|BBCUD4F_0|GNDO 0.07fF
C634 raven_soc_0|ram_rdata<23> raven_soc_0|ram_addr<0> 5.82fF
C635 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<15> 14.38fF
C636 BU_3VX2_71|Q raven_soc_0|flash_io3_oeb 0.02fF
C637 BU_3VX2_22|A BU_3VX2_20|Q 0.03fF
C638 BU_3VX2_0|A BU_3VX2_29|Q 0.02fF
C639 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<9> 0.02fF
C640 BU_3VX2_14|A raven_soc_0|flash_io3_do 0.01fF
C641 LS_3VX2_6|A LS_3VX2_16|A 0.01fF
C642 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<13> 0.02fF
C643 LOGIC0_3V_4|Q raven_padframe_0|ICF_1|PO 0.04fF
C644 raven_soc_0|gpio_out<2> BU_3VX2_25|Q 0.01fF
C645 BU_3VX2_7|A IN_3VX2_1|A 0.01fF
C646 BU_3VX2_8|A BU_3VX2_28|A 0.01fF
C647 LS_3VX2_3|Q BU_3VX2_18|A 0.01fF
C648 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<11> 1.31fF
C649 BU_3VX2_31|A BU_3VX2_0|Q 0.03fF
C650 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<5> 0.01fF
C651 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<7> 0.01fF
C652 raven_soc_0|gpio_outenb<4> BU_3VX2_71|Q 0.35fF
C653 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<13> 12.03fF
C654 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<8> 0.01fF
C655 BU_3VX2_73|Q LS_3VX2_17|A 0.01fF
C656 BU_3VX2_35|Q BU_3VX2_26|Q 0.01fF
C657 BU_3VX2_68|Q BU_3VX2_25|Q 0.05fF
C658 BU_3VX2_69|Q vdd 0.96fF
C659 BU_3VX2_56|Q vdd 2.00fF
C660 raven_soc_0|gpio_in<10> raven_padframe_0|BBCUD4F_10|PO 0.04fF
C661 BU_3VX2_16|A BU_3VX2_71|A 0.01fF
C662 BU_3VX2_1|A BU_3VX2_67|A 0.53fF
C663 BU_3VX2_71|A BU_3VX2_29|A 0.01fF
C664 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<3> 5.08fF
C665 BU_3VX2_31|A raven_soc_0|gpio_pulldown<0> 0.01fF
C666 BU_3VX2_5|A BU_3VX2_27|A 0.01fF
C667 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<9> 0.01fF
C668 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<16> 4.97fF
C669 raven_soc_0|ram_wdata<27> raven_soc_0|ram_wdata<31> 33.03fF
C670 raven_soc_0|ram_wdata<21> raven_soc_0|ram_addr<0> 0.01fF
C671 raven_soc_0|ram_wdata<25> raven_soc_0|ram_rdata<17> 0.01fF
C672 raven_soc_0|flash_io0_oeb vdd 2.65fF
C673 BU_3VX2_45|A BU_3VX2_43|A 1.80fF
C674 BU_3VX2_41|A LS_3VX2_27|Q 0.16fF
C675 BU_3VX2_46|A LS_3VX2_20|Q 0.35fF
C676 raven_soc_0|flash_io2_do BU_3VX2_28|Q 0.01fF
C677 raven_soc_0|flash_io2_oeb BU_3VX2_24|Q 0.01fF
C678 BU_3VX2_59|A BU_3VX2_60|Q 0.14fF
C679 raven_soc_0|gpio_out<15> BU_3VX2_27|Q 0.01fF
C680 AMUX4_3V_0|SEL[1] BU_3VX2_46|Q 26.00fF
C681 BU_3VX2_49|A BU_3VX2_49|Q 0.10fF
C682 BU_3VX2_46|Q BU_3VX2_51|Q 21.35fF
C683 BU_3VX2_37|A BU_3VX2_71|A 0.01fF
C684 raven_padframe_0|FILLER01F_0|VDDR raven_padframe_0|FILLER01F_0|GNDR 0.68fF
C685 raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# 0.22fF
C686 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<11> 0.01fF
C687 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<6> 0.01fF
C688 BU_3VX2_10|A raven_soc_0|flash_io2_do 0.03fF
C689 BU_3VX2_31|A BU_3VX2_30|Q 0.16fF
C690 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<15> 13.33fF
C691 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<5> 2.81fF
C692 raven_soc_0|gpio_pullup<9> BU_3VX2_40|Q 1.26fF
C693 LS_3VX2_3|A raven_soc_0|flash_io3_do 0.35fF
C694 raven_soc_0|gpio_pullup<8> raven_soc_0|ext_clk 0.01fF
C695 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<7> 2.63fF
C696 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<11> 0.02fF
C697 raven_soc_0|gpio_pullup<10> VDD3V3 0.07fF
C698 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<11> 5.03fF
C699 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<20> 5.26fF
C700 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<28> 7.17fF
C701 BU_3VX2_71|Q apllc03_1v8_0|CLK 32.34fF
C702 BU_3VX2_36|Q apllc03_1v8_0|CLK 1.00fF
C703 BU_3VX2_21|A BU_3VX2_20|Q 0.16fF
C704 LS_3VX2_11|A LS_3VX2_15|A 0.02fF
C705 IN_3VX2_1|Q BU_3VX2_62|Q 0.01fF
C706 BU_3VX2_40|A raven_soc_0|flash_io0_oeb 0.01fF
C707 BU_3VX2_0|A raven_soc_0|flash_io2_do 6.62fF
C708 BU_3VX2_18|A raven_soc_0|flash_io1_oeb 0.01fF
C709 LOGIC0_3V_4|Q raven_soc_0|gpio_in<14> 11.65fF
C710 BU_3VX2_31|A raven_soc_0|flash_io3_di 4.41fF
C711 BU_3VX2_13|A raven_soc_0|flash_io2_oeb 0.01fF
C712 VDD raven_padframe_0|FILLER50F_0|GNDO 0.07fF
C713 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<12> 1.89fF
C714 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<2> 10.66fF
C715 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pulldown<6> 4.99fF
C716 BU_3VX2_0|Q raven_soc_0|gpio_out<8> 0.50fF
C717 LS_3VX2_3|A raven_soc_0|gpio_out<14> 0.49fF
C718 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pulldown<7> 0.02fF
C719 BU_3VX2_0|Q BU_3VX2_3|Q 0.01fF
C720 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<9> 0.02fF
C721 BU_3VX2_33|A raven_soc_0|flash_io1_do 0.19fF
C722 LS_3VX2_13|A BU_3VX2_50|Q 5.09fF
C723 BU_3VX2_6|A BU_3VX2_13|A 1.60fF
C724 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<6> 0.01fF
C725 raven_soc_0|gpio_in<4> raven_soc_0|flash_io0_di 0.19fF
C726 AMUX2_3V_0|SEL LS_3VX2_27|A 14.29fF
C727 raven_soc_0|ram_rdata<12> vdd 0.59fF
C728 BU_3VX2_55|A BU_3VX2_54|Q 0.03fF
C729 LS_3VX2_22|A LS_3VX2_20|A 9.48fF
C730 acmpc01_3v3_0|IBN LS_3VX2_23|Q 6.15fF
C731 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<11> 0.01fF
C732 BU_3VX2_7|A BU_3VX2_25|A 0.01fF
C733 LS_3VX2_3|Q BU_3VX2_71|A 1.45fF
C734 BU_3VX2_8|A BU_3VX2_14|A 2.03fF
C735 LS_3VX2_10|A LS_3VX2_13|A 14.23fF
C736 VDD raven_soc_0|gpio_outenb<15> 0.20fF
C737 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<4> 4.07fF
C738 LS_3VX2_5|Q LS_3VX2_24|Q 0.01fF
C739 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_out<3> 1.86fF
C740 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<8> 0.01fF
C741 IN_3VX2_1|A raven_soc_0|gpio_pullup<15> 0.01fF
C742 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<6> 0.25fF
C743 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<10> 7.86fF
C744 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<7> 2.67fF
C745 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<5> 0.02fF
C746 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<11> 0.02fF
C747 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<13> 41.61fF
C748 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<15> 0.01fF
C749 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<11> 47.87fF
C750 BU_3VX2_0|Q raven_soc_0|gpio_out<6> 0.01fF
C751 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<7> 2.13fF
C752 raven_soc_0|gpio_out<1> BU_3VX2_28|Q 0.01fF
C753 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<21> 20.61fF
C754 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<10> 0.52fF
C755 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<7> 25.08fF
C756 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<22> 12.23fF
C757 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<20> 6.38fF
C758 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<23> 19.76fF
C759 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<9> 0.29fF
C760 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<30> 0.12fF
C761 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<24> 0.12fF
C762 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<14> 1.72fF
C763 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<4> 0.01fF
C764 raven_soc_0|flash_io3_do raven_soc_0|flash_io1_do 123.47fF
C765 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<15> 0.19fF
C766 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<25> 0.03fF
C767 BU_3VX2_14|Q BU_3VX2_9|Q 13.86fF
C768 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<17> 8.36fF
C769 BU_3VX2_70|Q BU_3VX2_69|Q 47.35fF
C770 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<14> 0.44fF
C771 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<12> 6.91fF
C772 BU_3VX2_15|Q BU_3VX2_14|Q 64.94fF
C773 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<2> 7.75fF
C774 BU_3VX2_32|Q BU_3VX2_5|Q 3.66fF
C775 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<1> 4.39fF
C776 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<13> 0.01fF
C777 BU_3VX2_16|Q BU_3VX2_3|Q 2.45fF
C778 BU_3VX2_35|Q BU_3VX2_11|Q 1.93fF
C779 BU_3VX2_26|Q BU_3VX2_23|Q 81.33fF
C780 vdd BU_3VX2_29|Q 4.35fF
C781 BU_3VX2_25|Q BU_3VX2_24|Q 349.59fF
C782 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<15> 30.91fF
C783 raven_padframe_0|aregc01_3v3_0|VDDR raven_padframe_0|aregc01_3v3_0|GNDO 0.10fF
C784 raven_padframe_0|aregc01_3v3_0|GNDR raven_padframe_0|aregc01_3v3_0|VDDO 0.07fF
C785 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<2> 7.11fF
C786 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<12> 0.01fF
C787 raven_soc_0|gpio_in<4> BU_3VX2_63|Q 0.01fF
C788 AMUX4_3V_1|AIN1 BU_3VX2_62|A 0.43fF
C789 BU_3VX2_19|A raven_soc_0|ext_clk 0.01fF
C790 VDD raven_padframe_0|GNDORPADF_1|VDDR 0.71fF
C791 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<23> 0.01fF
C792 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<31> 27.57fF
C793 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<1> 0.16fF
C794 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<13> 27.98fF
C795 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<29> 0.01fF
C796 VDD raven_soc_0|ser_tx 0.17fF
C797 VDD raven_padframe_0|FILLER01F_1|GNDR 0.16fF
C798 LS_3VX2_11|A AMUX4_3V_1|SEL[1] 14.85fF
C799 IN_3VX2_1|Q BU_3VX2_45|Q 1.03fF
C800 VDD raven_padframe_0|FILLER01F_0|GNDO 0.07fF
C801 BU_3VX2_26|A raven_soc_0|flash_io2_di 0.01fF
C802 VDD raven_padframe_0|aregc01_3v3_1|VDDR 0.54fF
C803 raven_soc_0|gpio_outenb<3> apllc03_1v8_0|CLK 0.01fF
C804 BU_3VX2_0|Q raven_soc_0|ram_rdata<18> 0.02fF
C805 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<8> 0.01fF
C806 raven_soc_0|gpio_in<2> BU_3VX2_29|Q 0.01fF
C807 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<12> 9.11fF
C808 BU_3VX2_63|Q raven_soc_0|gpio_in<7> 0.01fF
C809 BU_3VX2_27|A BU_3VX2_24|Q 0.02fF
C810 raven_soc_0|gpio_outenb<8> BU_3VX2_71|Q 0.01fF
C811 raven_padframe_0|BBCUD4F_6|VDDO raven_padframe_0|BBCUD4F_6|GNDO 2.28fF
C812 VDD raven_padframe_0|FILLER20F_8|VDDR 0.71fF
C813 LS_3VX2_11|A LS_3VX2_7|A 154.27fF
C814 LS_3VX2_6|Q LS_3VX2_5|Q 3.18fF
C815 BU_3VX2_63|A BU_3VX2_31|A 0.01fF
C816 LS_3VX2_10|A raven_soc_0|ser_rx 0.01fF
C817 raven_padframe_0|FILLER20F_0|VDDR raven_padframe_0|FILLER20F_0|GNDO 0.13fF
C818 raven_soc_0|gpio_pulldown<1> LS_3VX2_3|A 0.27fF
C819 BU_3VX2_22|A raven_soc_0|flash_io3_di 0.01fF
C820 AMUX4_3V_3|AOUT raven_soc_0|flash_io0_do 3.05fF
C821 raven_soc_0|gpio_pulldown<2> BU_3VX2_0|Q 0.01fF
C822 BU_3VX2_71|A raven_soc_0|flash_io1_oeb 0.01fF
C823 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<14> 0.46fF
C824 LOGIC0_3V_4|Q raven_soc_0|ser_tx 6.43fF
C825 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<3> 2.43fF
C826 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<6> 0.54fF
C827 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<13> 8.90fF
C828 BU_3VX2_11|A raven_soc_0|flash_io2_di 0.01fF
C829 raven_padframe_0|FILLER20F_5|VDDR raven_padframe_0|FILLER20F_5|GNDO 0.13fF
C830 BU_3VX2_24|A BU_3VX2_16|A 2.65fF
C831 BU_3VX2_24|A BU_3VX2_29|A 7.57fF
C832 raven_padframe_0|FILLER20F_8|VDDR LOGIC0_3V_4|Q 0.01fF
C833 LS_3VX2_8|Q LS_3VX2_5|Q 0.88fF
C834 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<5> 0.01fF
C835 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<2> 5.84fF
C836 BU_3VX2_13|A BU_3VX2_27|A 0.01fF
C837 BU_3VX2_24|A BU_3VX2_37|A 0.01fF
C838 raven_soc_0|ram_rdata<3> raven_soc_0|ram_addr<0> 0.04fF
C839 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<31> 0.02fF
C840 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<17> 7.72fF
C841 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<21> 0.01fF
C842 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<27> 0.01fF
C843 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<25> 0.01fF
C844 raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<22> 38.47fF
C845 raven_soc_0|ram_wdata<15> raven_soc_0|ram_rdata<15> 0.44fF
C846 raven_soc_0|ram_wdata<17> raven_soc_0|ram_rdata<1> 0.22fF
C847 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<17> 0.02fF
C848 raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<29> 11.52fF
C849 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<31> 21.44fF
C850 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<16> 7.62fF
C851 raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<13> 1.46fF
C852 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<27> 10.10fF
C853 raven_soc_0|flash_io2_do vdd 1.04fF
C854 BU_3VX2_50|A BU_3VX2_43|A 0.28fF
C855 BU_3VX2_51|A LS_3VX2_21|Q 0.11fF
C856 BU_3VX2_59|A BU_3VX2_62|Q 0.02fF
C857 raven_soc_0|gpio_in<11> BU_3VX2_29|Q 0.01fF
C858 raven_soc_0|gpio_out<15> BU_3VX2_25|Q 0.01fF
C859 BU_3VX2_46|Q BU_3VX2_49|Q 32.73fF
C860 BU_3VX2_43|Q BU_3VX2_72|Q 0.29fF
C861 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<8> 0.01fF
C862 raven_padframe_0|VDDPADF_1|GNDR raven_padframe_0|VDDPADF_1|GNDO 0.81fF
C863 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<2> 0.74fF
C864 raven_padframe_0|axtoc02_3v3_0|m4_55000_31172# raven_padframe_0|axtoc02_3v3_0|m4_55000_30653# 0.17fF
C865 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<11> 0.01fF
C866 BU_3VX2_63|Q raven_soc_0|gpio_out<7> 0.01fF
C867 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<5> 0.01fF
C868 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<5> 0.01fF
C869 BU_3VX2_1|A BU_3VX2_33|Q 0.16fF
C870 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<14> 31.98fF
C871 raven_soc_0|gpio_pulldown<9> BU_3VX2_40|Q 0.17fF
C872 raven_soc_0|gpio_pulldown<4> VDD3V3 0.09fF
C873 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<12> 8.55fF
C874 BU_3VX2_1|Q raven_soc_0|flash_clk 0.63fF
C875 BU_3VX2_70|Q BU_3VX2_29|Q 0.65fF
C876 BU_3VX2_4|Q BU_3VX2_26|Q 0.02fF
C877 BU_3VX2_32|Q BU_3VX2_28|Q 0.45fF
C878 LS_3VX2_22|A BU_3VX2_47|Q 5.17fF
C879 raven_soc_0|gpio_out<10> BU_3VX2_27|Q 0.01fF
C880 BU_3VX2_11|Q BU_3VX2_23|Q 3.05fF
C881 raven_soc_0|gpio_outenb<13> BU_3VX2_23|Q 0.01fF
C882 raven_soc_0|gpio_pullup<14> apllc03_1v8_0|CLK 0.01fF
C883 raven_soc_0|gpio_outenb<9> BU_3VX2_29|Q 0.01fF
C884 BU_3VX2_23|A BU_3VX2_22|Q 0.16fF
C885 BU_3VX2_8|A raven_soc_0|flash_io1_do 0.01fF
C886 BU_3VX2_40|A raven_soc_0|flash_io2_do 0.01fF
C887 raven_padframe_0|BBC4F_2|VDDR raven_padframe_0|BBC4F_2|VDDO 0.06fF
C888 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<13> 0.73fF
C889 LS_3VX2_8|A AMUX4_3V_4|AIN2 0.63fF
C890 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pulldown<7> 0.01fF
C891 LS_3VX2_7|A LS_3VX2_21|A 7.82fF
C892 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<7> 0.36fF
C893 BU_3VX2_0|Q raven_soc_0|gpio_pulldown<6> 0.01fF
C894 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<6> 0.01fF
C895 BU_3VX2_47|A BU_3VX2_46|A 2.92fF
C896 BU_3VX2_7|A BU_3VX2_4|A 4.64fF
C897 BU_3VX2_21|A raven_soc_0|flash_io3_di 0.11fF
C898 BU_3VX2_17|A raven_soc_0|flash_io0_do 0.01fF
C899 raven_soc_0|gpio_out<0> apllc03_1v8_0|B_CP 0.01fF
C900 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<8> 0.33fF
C901 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<6> 2.86fF
C902 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<6> 0.60fF
C903 raven_padframe_0|ICF_0|VDDR raven_padframe_0|ICF_0|GNDO 0.13fF
C904 LS_3VX2_13|A raven_soc_0|ser_tx 0.01fF
C905 raven_soc_0|gpio_out<11> BU_3VX2_28|Q 0.01fF
C906 raven_soc_0|gpio_out<9> BU_3VX2_27|Q 0.01fF
C907 BU_3VX2_24|A LS_3VX2_3|Q 0.01fF
C908 BU_3VX2_73|Q BU_3VX2_42|Q 24.77fF
C909 BU_3VX2_55|A BU_3VX2_56|Q 0.15fF
C910 BU_3VX2_22|A BU_3VX2_63|A 0.02fF
C911 VDD3V3 raven_padframe_0|VDDORPADF_3|GNDR 0.78fF
C912 raven_soc_0|gpio_out<0> LS_3VX2_3|A 0.13fF
C913 BU_3VX2_16|A BU_3VX2_29|A 1.59fF
C914 LS_3VX2_24|A LS_3VX2_13|A 23.27fF
C915 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<11> 0.80fF
C916 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<12> 0.03fF
C917 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<10> 7.86fF
C918 LS_3VX2_3|A raven_soc_0|gpio_out<12> 0.01fF
C919 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<14> 0.02fF
C920 BU_3VX2_0|Q raven_soc_0|gpio_outenb<11> 0.01fF
C921 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<7> 2.63fF
C922 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<15> 15.53fF
C923 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<11> 10.57fF
C924 raven_soc_0|gpio_out<1> vdd 0.50fF
C925 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<10> 0.01fF
C926 AMUX4_3V_3|SEL[1] BU_3VX2_67|Q 0.20fF
C927 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<25> 32.23fF
C928 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<8> 0.42fF
C929 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<8> 0.11fF
C930 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<4> 0.10fF
C931 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<2> 0.07fF
C932 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<12> 3.91fF
C933 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<1> 0.01fF
C934 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<21> 0.05fF
C935 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<7> 0.47fF
C936 BU_3VX2_40|Q raven_soc_0|flash_io0_di 24.22fF
C937 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<5> 0.01fF
C938 BU_3VX2_14|Q BU_3VX2_64|Q 37.33fF
C939 raven_soc_0|flash_io2_di VDD3V3 9.21fF
C940 VDD3V3 AMUX4_3V_0|AOUT 6.55fF
C941 BU_3VX2_50|Q BU_3VX2_72|Q 2.61fF
C942 acsoc02_3v3_0|CS_4U aopac01_3v3_0|IB 0.49fF
C943 BU_3VX2_37|A BU_3VX2_29|A 0.01fF
C944 BU_3VX2_72|A IN_3VX2_1|A 0.01fF
C945 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<7> 0.29fF
C946 BU_3VX2_33|A raven_soc_0|flash_csb 0.01fF
C947 AMUX4_3V_1|AIN1 BU_3VX2_55|A 0.02fF
C948 BU_3VX2_12|A BU_3VX2_12|Q 0.08fF
C949 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<23> 14.95fF
C950 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<10> 0.12fF
C951 BU_3VX2_71|Q raven_soc_0|gpio_in<15> 0.02fF
C952 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<20> 0.01fF
C953 BU_3VX2_1|Q BU_3VX2_61|Q 0.56fF
C954 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<19> 1.04fF
C955 raven_soc_0|ram_wdata<24> vdd 1.07fF
C956 BU_3VX2_59|Q BU_3VX2_53|Q 23.60fF
C957 raven_soc_0|ram_wdata<23> apllc03_1v8_0|CLK 0.01fF
C958 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<2> 9.22fF
C959 LS_3VX2_9|A BU_3VX2_54|Q 16.32fF
C960 IN_3VX2_1|Q AMUX4_3V_4|AIN3 6.59fF
C961 AMUX4_3V_0|AIN1 BU_3VX2_44|A 0.02fF
C962 BU_3VX2_12|A raven_soc_0|flash_io0_do 0.01fF
C963 BU_3VX2_69|A BU_3VX2_69|Q 0.08fF
C964 BU_3VX2_63|Q BU_3VX2_40|Q 113.39fF
C965 raven_soc_0|gpio_pulldown<11> VDD3V3 0.07fF
C966 raven_soc_0|ser_rx raven_soc_0|ser_tx 485.01fF
C967 BU_3VX2_31|A BU_3VX2_26|Q 31.55fF
C968 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<6> 67.13fF
C969 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<10> 0.12fF
C970 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<24> 0.31fF
C971 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<31> 14.09fF
C972 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_outenb<8> 0.74fF
C973 BU_3VX2_11|Q BU_3VX2_4|Q 7.23fF
C974 raven_padframe_0|FILLER10F_1|VDDR raven_padframe_0|FILLER10F_1|VDDO 0.06fF
C975 markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# markings_0|manufacturer_0|_alphabet_E_1|m2_0_0# 0.01fF
C976 BU_3VX2_24|A raven_soc_0|flash_io1_oeb 3.27fF
C977 BU_3VX2_38|A BU_3VX2_26|A 0.37fF
C978 LS_3VX2_24|A raven_soc_0|ser_rx 0.01fF
C979 BU_3VX2_3|A raven_soc_0|flash_io0_di 0.01fF
C980 BU_3VX2_15|A raven_soc_0|flash_io0_di 0.01fF
C981 raven_soc_0|gpio_pullup<2> BU_3VX2_29|Q 0.01fF
C982 raven_soc_0|gpio_in<3> raven_soc_0|flash_io2_oeb 5.25fF
C983 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<7> 1.89fF
C984 raven_soc_0|gpio_in<0> raven_soc_0|flash_io3_do 0.17fF
C985 raven_soc_0|flash_csb raven_soc_0|flash_io3_do 14.60fF
C986 raven_soc_0|flash_csb AMUX4_3V_4|AIN3 7.87fF
C987 BU_3VX2_21|A BU_3VX2_63|A 0.01fF
C988 BU_3VX2_16|A LS_3VX2_3|Q 0.01fF
C989 BU_3VX2_38|A LOGIC0_3V_3|Q 0.01fF
C990 BU_3VX2_38|A BU_3VX2_11|A 1.92fF
C991 LS_3VX2_3|Q BU_3VX2_29|A 0.01fF
C992 LS_3VX2_12|Q LS_3VX2_24|Q 0.01fF
C993 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<2> 14.70fF
C994 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<14> 0.09fF
C995 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<11> 0.16fF
C996 raven_soc_0|gpio_out<13> BU_3VX2_71|Q 0.01fF
C997 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<5> 14.65fF
C998 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<8> 0.01fF
C999 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<27> 38.99fF
C1000 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<13> 0.16fF
C1001 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<31> 40.44fF
C1002 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<29> 4.14fF
C1003 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<26> 0.01fF
C1004 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<1> 0.01fF
C1005 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<17> 0.01fF
C1006 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<19> 0.01fF
C1007 BU_3VX2_1|Q BU_3VX2_33|Q 51.67fF
C1008 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<22> 5.72fF
C1009 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<19> 13.75fF
C1010 raven_soc_0|ram_wdata<8> raven_soc_0|ram_rdata<1> 0.11fF
C1011 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<13> 0.01fF
C1012 raven_soc_0|gpio_in<9> apllc03_1v8_0|CLK 0.02fF
C1013 comp_inp AMUX4_3V_4|AIN2 130.33fF
C1014 raven_soc_0|ext_clk BU_3VX2_27|Q 0.01fF
C1015 raven_soc_0|gpio_in<12> BU_3VX2_28|Q 0.01fF
C1016 BU_3VX2_37|A LS_3VX2_3|Q 0.01fF
C1017 raven_padframe_0|GNDORPADF_2|VDDR raven_padframe_0|GNDORPADF_2|VDDO 0.06fF
C1018 raven_padframe_0|aregc01_3v3_1|m4_92500_30653# raven_padframe_0|aregc01_3v3_1|m4_92500_29333# 0.02fF
C1019 raven_padframe_0|aregc01_3v3_1|m4_0_29333# raven_padframe_0|aregc01_3v3_1|m4_0_22024# 0.01fF
C1020 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<3> 3.29fF
C1021 raven_padframe_0|axtoc02_3v3_0|m4_0_29057# raven_padframe_0|axtoc02_3v3_0|m4_0_28769# 0.22fF
C1022 BU_3VX2_63|Q raven_soc_0|gpio_outenb<7> 0.01fF
C1023 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<11> 0.01fF
C1024 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<7> 11.71fF
C1025 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<6> 0.01fF
C1026 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<9> 0.03fF
C1027 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<8> 0.07fF
C1028 LS_3VX2_3|A raven_soc_0|gpio_pullup<5> 0.08fF
C1029 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<12> 172.99fF
C1030 raven_soc_0|gpio_out<10> BU_3VX2_25|Q 0.01fF
C1031 raven_soc_0|gpio_pullup<13> BU_3VX2_23|Q 0.01fF
C1032 BU_3VX2_32|Q vdd 1.58fF
C1033 BU_3VX2_3|Q BU_3VX2_26|Q 0.01fF
C1034 BU_3VX2_37|Q BU_3VX2_24|Q 0.01fF
C1035 BU_3VX2_20|A raven_soc_0|flash_io3_do 0.01fF
C1036 BU_3VX2_7|A raven_soc_0|flash_io0_oeb 0.01fF
C1037 LS_3VX2_10|A AMUX4_3V_1|SEL[0] 18.66fF
C1038 raven_padframe_0|BBC4F_1|VDDR raven_padframe_0|BBC4F_1|GNDR 0.68fF
C1039 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<13> 0.01fF
C1040 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<7> 1.03fF
C1041 LS_3VX2_7|A LS_3VX2_27|A 8.36fF
C1042 raven_soc_0|gpio_out<2> BU_3VX2_40|Q 0.02fF
C1043 raven_padframe_0|BBCUD4F_10|VDDR raven_padframe_0|BBCUD4F_10|GNDO 0.13fF
C1044 BU_3VX2_26|A BU_3VX2_23|Q 0.02fF
C1045 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<20> 9.96fF
C1046 BU_3VX2_48|A adc0_data<5> 0.04fF
C1047 raven_padframe_0|APR00DF_4|VDDR raven_padframe_0|APR00DF_4|GNDO 0.13fF
C1048 LS_3VX2_12|Q LS_3VX2_6|Q 2.51fF
C1049 BU_3VX2_23|A raven_soc_0|flash_io3_oeb 0.01fF
C1050 BU_3VX2_37|A BU_3VX2_38|Q 0.16fF
C1051 BU_3VX2_25|A BU_3VX2_22|Q 0.02fF
C1052 BU_3VX2_16|A raven_soc_0|flash_io1_oeb 0.01fF
C1053 IN_3VX2_1|Q LS_3VX2_21|A 0.01fF
C1054 BU_3VX2_17|A raven_soc_0|flash_io1_di 0.08fF
C1055 BU_3VX2_31|A raven_soc_0|gpio_outenb<13> 0.01fF
C1056 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<15> 0.12fF
C1057 BU_3VX2_29|A raven_soc_0|flash_io1_oeb 8.08fF
C1058 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<3> 1.66fF
C1059 VDD raven_padframe_0|APR00DF_4|GNDR 0.16fF
C1060 raven_soc_0|gpio_out<11> vdd 0.19fF
C1061 raven_soc_0|gpio_outenb<10> BU_3VX2_27|Q 0.01fF
C1062 AMUX2_3V_0|SEL BU_3VX2_53|Q 0.01fF
C1063 raven_soc_0|gpio_outenb<14> BU_3VX2_29|Q 0.01fF
C1064 raven_soc_0|gpio_out<9> BU_3VX2_25|Q 0.01fF
C1065 BU_3VX2_23|A BU_3VX2_2|A 0.01fF
C1066 LS_3VX2_9|A LS_3VX2_14|A 9.88fF
C1067 LS_3VX2_8|Q LS_3VX2_12|Q 16.47fF
C1068 BU_3VX2_32|A BU_3VX2_65|A 0.53fF
C1069 LS_3VX2_19|Q acsoc02_3v3_0|CS_8U 0.06fF
C1070 LS_3VX2_5|Q LS_3VX2_14|Q 1.03fF
C1071 LS_3VX2_10|Q LS_3VX2_7|A 0.18fF
C1072 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<5> 2.97fF
C1073 BU_3VX2_37|A raven_soc_0|flash_io1_oeb 0.01fF
C1074 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<9> 122.66fF
C1075 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<8> 0.03fF
C1076 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<4> 0.14fF
C1077 LS_3VX2_3|A raven_soc_0|gpio_outenb<12> 0.01fF
C1078 BU_3VX2_0|Q raven_soc_0|gpio_pullup<11> 0.01fF
C1079 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<15> 0.02fF
C1080 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<5> 5.77fF
C1081 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<8> 0.31fF
C1082 LOGIC0_3V_1|Q LOGIC1_3V_0|Q 2.88fF
C1083 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<0> 0.43fF
C1084 raven_soc_0|gpio_in<7> raven_soc_0|gpio_out<15> 0.24fF
C1085 AMUX4_3V_3|SEL[1] BU_3VX2_65|Q 0.18fF
C1086 raven_soc_0|ext_clk raven_soc_0|flash_io2_oeb 20.57fF
C1087 raven_soc_0|irq_pin BU_3VX2_52|Q 0.01fF
C1088 AMUX4_3V_4|AIN2 vdd 8.34fF
C1089 BU_3VX2_48|Q BU_3VX2_72|Q 1.97fF
C1090 LS_3VX2_20|A BU_3VX2_45|Q 11.20fF
C1091 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<2> 17.39fF
C1092 BU_3VX2_3|A BU_3VX2_5|A 7.43fF
C1093 VDD LOGIC0_3V_4|Q 1.39fF
C1094 BU_3VX2_5|A BU_3VX2_15|A 1.06fF
C1095 BU_3VX2_8|A raven_soc_0|flash_csb 0.01fF
C1096 raven_padframe_0|BBCUD4F_5|VDDO raven_padframe_0|BBCUD4F_5|GNDO 2.28fF
C1097 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_in<0> 11.29fF
C1098 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<13> 0.01fF
C1099 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<5> 6.64fF
C1100 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<11> 2.80fF
C1101 raven_padframe_0|aregc01_3v3_0|m4_92500_30133# raven_padframe_0|aregc01_3v3_0|m4_92500_29333# 0.09fF
C1102 raven_padframe_0|aregc01_3v3_0|m4_92500_30653# raven_padframe_0|aregc01_3v3_0|m4_92500_29057# 0.01fF
C1103 raven_padframe_0|aregc01_3v3_0|m4_0_28769# raven_padframe_0|aregc01_3v3_0|m4_0_22024# 0.03fF
C1104 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<7> 0.01fF
C1105 markings_0|efabless_logo_0|m2_4800_n4350# markings_0|efabless_logo_0|m2_3000_n6450# 0.41fF
C1106 BU_3VX2_6|A raven_soc_0|ext_clk 0.04fF
C1107 BU_3VX2_38|A VDD3V3 0.31fF
C1108 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<25> 56.62fF
C1109 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<0> 10.65fF
C1110 BU_3VX2_71|Q raven_soc_0|gpio_in<14> 0.02fF
C1111 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<15> 0.04fF
C1112 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<7> 3.80fF
C1113 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<13> 44.27fF
C1114 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<17> 0.05fF
C1115 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<9> 6.87fF
C1116 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<2> 1.90fF
C1117 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<15> 50.05fF
C1118 BU_3VX2_61|Q BU_3VX2_53|Q 15.90fF
C1119 raven_soc_0|ram_rdata<8> vdd 0.30fF
C1120 LS_3VX2_18|A apllc03_1v8_0|CLK 0.59fF
C1121 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<8> 0.11fF
C1122 LS_3VX2_9|A BU_3VX2_56|Q 10.97fF
C1123 LS_3VX2_10|A LS_3VX2_17|A 0.01fF
C1124 BU_3VX2_12|A raven_soc_0|flash_io1_di 0.01fF
C1125 IN_3VX2_1|A BU_3VX2_31|Q 0.03fF
C1126 adc_low raven_soc_0|irq_pin 0.05fF
C1127 raven_soc_0|gpio_pullup<0> apllc03_1v8_0|CLK 0.02fF
C1128 raven_soc_0|gpio_pulldown<2> BU_3VX2_26|Q 0.01fF
C1129 raven_soc_0|gpio_out<8> raven_soc_0|gpio_outenb<13> 0.51fF
C1130 raven_soc_0|gpio_pullup<6> BU_3VX2_71|Q 0.10fF
C1131 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<10> 4.78fF
C1132 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<6> 18.93fF
C1133 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<24> 0.70fF
C1134 raven_soc_0|ram_addr<3> raven_soc_0|ram_addr<2> 94.97fF
C1135 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<9> 2.68fF
C1136 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<7> 0.05fF
C1137 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<31> 0.02fF
C1138 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<20> 0.01fF
C1139 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<6> 0.01fF
C1140 BU_3VX2_3|Q BU_3VX2_11|Q 17.40fF
C1141 BU_3VX2_70|Q BU_3VX2_32|Q 0.45fF
C1142 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<2> 5.92fF
C1143 markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# 1.06fF
C1144 markings_0|product_name_0|_alphabet_V_1|m2_0_560# markings_0|product_name_0|_alphabet_N_0|m2_0_0# 0.09fF
C1145 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<10> 3.61fF
C1146 AMUX4_3V_3|AOUT comp_inp 0.36fF
C1147 LS_3VX2_3|Q raven_soc_0|flash_io1_oeb 0.01fF
C1148 IN_3VX2_1|A raven_soc_0|flash_io3_oeb 6.87fF
C1149 LS_3VX2_6|A LS_3VX2_19|A 0.01fF
C1150 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<11> 50.22fF
C1151 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<10> 9.74fF
C1152 LS_3VX2_6|A BU_3VX2_52|Q 12.79fF
C1153 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<15> 0.02fF
C1154 BU_3VX2_0|Q raven_soc_0|ram_rdata<20> 0.02fF
C1155 BU_3VX2_8|A BU_3VX2_20|A 0.98fF
C1156 BU_3VX2_10|A BU_3VX2_17|A 1.83fF
C1157 BU_3VX2_2|A IN_3VX2_1|A 0.01fF
C1158 raven_padframe_0|ICFC_1|VDD3 BU_3VX2_33|A 0.01fF
C1159 AMUX4_3V_0|AIN1 BU_3VX2_48|A 0.02fF
C1160 BU_3VX2_71|A BU_3VX2_71|Q 0.09fF
C1161 LOGIC0_3V_4|Q raven_soc_0|flash_io1_oeb 0.01fF
C1162 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<5> 0.50fF
C1163 raven_soc_0|gpio_outenb<15> BU_3VX2_71|Q 0.01fF
C1164 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pullup<14> 12.44fF
C1165 raven_soc_0|gpio_out<11> raven_soc_0|gpio_outenb<9> 6.25fF
C1166 raven_soc_0|gpio_out<6> raven_soc_0|gpio_outenb<13> 0.01fF
C1167 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<29> 1.38fF
C1168 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<27> 164.47fF
C1169 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<1> 0.01fF
C1170 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<7> 0.01fF
C1171 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<6> 0.01fF
C1172 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<5> 0.01fF
C1173 BU_3VX2_12|Q BU_3VX2_2|Q 6.70fF
C1174 BU_3VX2_13|Q BU_3VX2_22|Q 15.41fF
C1175 BU_3VX2_66|Q BU_3VX2_9|Q 1.33fF
C1176 BU_3VX2_6|Q BU_3VX2_8|Q 24.92fF
C1177 BU_3VX2_12|Q BU_3VX2_10|Q 23.68fF
C1178 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<26> 27.59fF
C1179 BU_3VX2_15|Q BU_3VX2_20|Q 7.08fF
C1180 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<27> 0.39fF
C1181 BU_3VX2_21|Q BU_3VX2_7|Q 0.12fF
C1182 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<13> 0.03fF
C1183 BU_3VX2_38|Q BU_3VX2_67|Q 0.01fF
C1184 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<19> 8.90fF
C1185 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<22> 4.92fF
C1186 BU_3VX2_7|Q BU_3VX2_8|Q 68.71fF
C1187 BU_3VX2_9|Q BU_3VX2_20|Q 2.87fF
C1188 raven_soc_0|gpio_in<12> vdd 2.52fF
C1189 VDD3V3 LS_3VX2_16|A 0.47fF
C1190 BU_3VX2_58|A vdd 0.29fF
C1191 raven_soc_0|ext_clk BU_3VX2_25|Q 0.01fF
C1192 VDD3V3 BU_3VX2_23|Q 0.82fF
C1193 BU_3VX2_40|Q BU_3VX2_24|Q 0.01fF
C1194 VDD raven_padframe_0|BT4F_1|VDDR 0.71fF
C1195 raven_padframe_0|FILLER50F_2|GNDR raven_padframe_0|FILLER50F_2|GNDO 0.81fF
C1196 VDD raven_padframe_0|BBCUD4F_2|VDDR 0.71fF
C1197 raven_padframe_0|FILLER20F_7|GNDR raven_padframe_0|FILLER20F_7|GNDO 0.81fF
C1198 BU_3VX2_0|A BU_3VX2_17|A 0.11fF
C1199 raven_padframe_0|aregc01_3v3_1|m4_0_30133# raven_padframe_0|aregc01_3v3_1|m4_0_29057# 0.01fF
C1200 raven_padframe_0|APR00DF_2|VDDR raven_padframe_0|APR00DF_2|VDDO 0.06fF
C1201 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<5> 0.65fF
C1202 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<4> 0.01fF
C1203 BU_3VX2_63|Q raven_soc_0|gpio_pullup<9> 0.01fF
C1204 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<8> 0.01fF
C1205 raven_soc_0|gpio_pulldown<8> BU_3VX2_0|Q 0.01fF
C1206 raven_soc_0|gpio_out<4> VDD3V3 0.24fF
C1207 raven_soc_0|irq_pin BU_3VX2_58|Q 0.01fF
C1208 raven_soc_0|gpio_pulldown<7> BU_3VX2_28|Q 0.01fF
C1209 raven_soc_0|ram_rdata<16> vdd 0.30fF
C1210 raven_soc_0|ram_wdata<31> apllc03_1v8_0|CLK 0.01fF
C1211 raven_padframe_0|BT4F_1|VDDR LOGIC0_3V_4|Q 0.01fF
C1212 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<0> 57.49fF
C1213 raven_padframe_0|BBCUD4F_2|VDDR LOGIC0_3V_4|Q 0.01fF
C1214 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<8> 0.26fF
C1215 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<12> 0.37fF
C1216 raven_padframe_0|VDDPADFC_0|VDDR VDD3V3 0.71fF
C1217 BU_3VX2_7|A raven_soc_0|flash_io2_do 0.01fF
C1218 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<12> 3.06fF
C1219 LS_3VX2_24|A AMUX4_3V_1|SEL[0] 0.12fF
C1220 BU_3VX2_31|A raven_soc_0|gpio_in<8> 0.01fF
C1221 VDD raven_padframe_0|BBCUD4F_10|GNDR 0.16fF
C1222 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<7> 1.28fF
C1223 BU_3VX2_0|Q raven_soc_0|ram_wdata<17> 0.02fF
C1224 BU_3VX2_27|A raven_soc_0|ext_clk 0.01fF
C1225 raven_soc_0|flash_io0_di raven_soc_0|ram_rdata<11> 14.79fF
C1226 raven_soc_0|ram_rdata<31> raven_soc_0|ram_addr<0> 92.58fF
C1227 raven_soc_0|flash_io0_do raven_soc_0|flash_clk 50.14fF
C1228 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<16> 2.64fF
C1229 BU_3VX2_45|A BU_3VX2_45|Q 0.10fF
C1230 BU_3VX2_45|Q BU_3VX2_47|Q 45.51fF
C1231 raven_padframe_0|BBCUD4F_4|GNDR raven_padframe_0|BBCUD4F_4|VDDO 0.09fF
C1232 raven_padframe_0|FILLER10F_0|GNDR raven_padframe_0|FILLER10F_0|GNDO 0.81fF
C1233 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<14> 0.51fF
C1234 BU_3VX2_10|A BU_3VX2_12|A 7.93fF
C1235 BU_3VX2_68|A BU_3VX2_70|A 8.53fF
C1236 BU_3VX2_9|A raven_soc_0|flash_io0_do 0.01fF
C1237 BU_3VX2_19|A raven_soc_0|flash_io2_di 0.01fF
C1238 AMUX4_3V_3|AOUT vdd 0.41fF
C1239 IN_3VX2_1|Q LS_3VX2_27|A 0.01fF
C1240 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<8> 0.19fF
C1241 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<6> 0.02fF
C1242 BU_3VX2_31|A raven_soc_0|gpio_pullup<13> 0.01fF
C1243 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<6> 9.30fF
C1244 IN_3VX2_1|A apllc03_1v8_0|CLK 3.51fF
C1245 VDD raven_padframe_0|FILLER20F_2|GNDO 0.07fF
C1246 raven_padframe_0|BBCUD4F_12|VDDR raven_padframe_0|BBCUD4F_12|VDDO 0.06fF
C1247 VDD raven_padframe_0|FILLER20F_3|GNDR 0.16fF
C1248 raven_soc_0|gpio_outenb<10> BU_3VX2_25|Q 0.01fF
C1249 raven_soc_0|gpio_pullup<15> BU_3VX2_29|Q 0.01fF
C1250 raven_soc_0|gpio_pullup<10> BU_3VX2_27|Q 0.01fF
C1251 raven_soc_0|gpio_outenb<11> BU_3VX2_26|Q 0.01fF
C1252 LS_3VX2_7|Q LS_3VX2_5|Q 1.38fF
C1253 VDD raven_soc_0|ser_rx 0.17fF
C1254 BU_3VX2_0|A BU_3VX2_12|A 0.01fF
C1255 BU_3VX2_31|A BU_3VX2_26|A 6.74fF
C1256 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<6> 0.83fF
C1257 LS_3VX2_3|A raven_soc_0|gpio_pullup<12> 0.01fF
C1258 BU_3VX2_25|A raven_soc_0|flash_io3_oeb 2.71fF
C1259 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<4> 0.01fF
C1260 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<10> 0.34fF
C1261 LS_3VX2_6|A BU_3VX2_58|Q 7.40fF
C1262 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<10> 3.90fF
C1263 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<15> 1.25fF
C1264 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<11> 21.38fF
C1265 raven_soc_0|gpio_in<7> raven_soc_0|gpio_in<6> 24.61fF
C1266 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<10> 0.02fF
C1267 BU_3VX2_40|Q raven_soc_0|gpio_out<15> 0.01fF
C1268 BU_3VX2_61|A LS_3VX2_15|Q 2.84fF
C1269 BU_3VX2_58|A BU_3VX2_62|A 0.24fF
C1270 BU_3VX2_59|A LS_3VX2_17|Q 0.23fF
C1271 BU_3VX2_60|A LS_3VX2_16|Q 0.45fF
C1272 AMUX4_3V_1|AOUT AMUX4_3V_4|AIN3 1.22fF
C1273 BU_3VX2_42|Q BU_3VX2_43|Q 63.55fF
C1274 BU_3VX2_2|A BU_3VX2_25|A 0.01fF
C1275 BU_3VX2_3|A BU_3VX2_13|A 0.99fF
C1276 raven_padframe_0|APR00DF_5|VDDR raven_padframe_0|APR00DF_5|GNDO 0.13fF
C1277 BU_3VX2_15|A BU_3VX2_13|A 12.14fF
C1278 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<13> 0.01fF
C1279 raven_padframe_0|FILLER20F_4|VDDR raven_padframe_0|FILLER20F_4|VDDO 0.06fF
C1280 LOGIC0_3V_4|Q raven_soc_0|ser_rx 7.11fF
C1281 BU_3VX2_31|A BU_3VX2_11|A 0.01fF
C1282 raven_padframe_0|aregc01_3v3_0|m4_0_29333# raven_padframe_0|aregc01_3v3_0|m4_0_29057# 0.11fF
C1283 raven_padframe_0|aregc01_3v3_0|m4_0_30133# raven_padframe_0|aregc01_3v3_0|m4_0_28769# 0.01fF
C1284 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<15> 0.29fF
C1285 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<7> 0.52fF
C1286 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<9> 0.01fF
C1287 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<19> 0.25fF
C1288 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<7> 2.55fF
C1289 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<8> 23.83fF
C1290 raven_soc_0|gpio_in<5> BU_3VX2_40|Q 0.01fF
C1291 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<11> 0.01fF
C1292 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<12> 0.02fF
C1293 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<14> 79.28fF
C1294 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<0> 4.01fF
C1295 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<2> 0.01fF
C1296 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<1> 0.79fF
C1297 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<12> 1.29fF
C1298 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<8> 0.04fF
C1299 raven_soc_0|ram_rdata<22> vdd 0.75fF
C1300 raven_soc_0|ser_tx LS_3VX2_17|A 44.96fF
C1301 LS_3VX2_15|A BU_3VX2_53|Q 10.63fF
C1302 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<1> 0.01fF
C1303 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<3> 5.71fF
C1304 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<9> 0.88fF
C1305 LS_3VX2_24|A LS_3VX2_17|A 0.01fF
C1306 BU_3VX2_0|Q BU_3VX2_15|Q 0.01fF
C1307 BU_3VX2_0|Q BU_3VX2_9|Q 0.01fF
C1308 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_pullup<14> 0.58fF
C1309 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_out<8> 0.02fF
C1310 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_outenb<13> 0.02fF
C1311 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<23> 3.20fF
C1312 AMUX4_3V_3|SEL[1] BU_3VX2_36|Q 0.16fF
C1313 raven_soc_0|ram_rdata<21> raven_soc_0|ram_addr<4> 0.13fF
C1314 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<9> 21.44fF
C1315 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<30> 0.02fF
C1316 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<8> 0.01fF
C1317 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<20> 0.01fF
C1318 raven_soc_0|ram_rdata<18> raven_soc_0|ram_addr<3> 0.01fF
C1319 raven_padframe_0|ICFC_2|VDDO raven_padframe_0|ICFC_2|GNDO 2.28fF
C1320 markings_0|manufacturer_0|_alphabet_E_2|m2_0_0# markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# 0.12fF
C1321 raven_soc_0|gpio_in<1> raven_soc_0|flash_io3_do 0.38fF
C1322 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<13> 4.01fF
C1323 BU_3VX2_17|A vdd 0.06fF
C1324 LS_3VX2_6|A LS_3VX2_22|A 11.00fF
C1325 BU_3VX2_28|A raven_soc_0|flash_io0_do 4.57fF
C1326 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<5> 0.01fF
C1327 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<9> 1.02fF
C1328 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<10> 8.04fF
C1329 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<7> 3.96fF
C1330 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<8> 1.33fF
C1331 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<13> 14.86fF
C1332 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<7> 0.89fF
C1333 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<6> 5.66fF
C1334 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<15> 0.02fF
C1335 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<14> 0.36fF
C1336 LS_3VX2_12|Q LS_3VX2_14|Q 0.35fF
C1337 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_outenb<1> 40.82fF
C1338 AMUX4_3V_0|AIN1 AMUX4_3V_0|AOUT 0.90fF
C1339 IN_3VX2_1|A raven_soc_0|gpio_outenb<8> 0.01fF
C1340 LS_3VX2_8|A BU_3VX2_59|Q 0.46fF
C1341 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<5> 0.06fF
C1342 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<8> 0.93fF
C1343 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<10> 1.13fF
C1344 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<13> 11.86fF
C1345 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<14> 0.72fF
C1346 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pullup<14> 84.34fF
C1347 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pullup<13> 0.01fF
C1348 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<27> 0.43fF
C1349 BU_3VX2_19|Q BU_3VX2_6|Q 3.64fF
C1350 BU_3VX2_16|Q BU_3VX2_15|Q 69.72fF
C1351 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<2> 0.31fF
C1352 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<30> 68.34fF
C1353 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<25> 0.03fF
C1354 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<29> 0.54fF
C1355 BU_3VX2_2|Q BU_3VX2_5|Q 17.42fF
C1356 BU_3VX2_66|Q BU_3VX2_64|Q 16.43fF
C1357 BU_3VX2_19|Q BU_3VX2_7|Q 4.46fF
C1358 BU_3VX2_6|Q BU_3VX2_18|Q 3.02fF
C1359 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<2> 0.23fF
C1360 BU_3VX2_13|Q BU_3VX2_31|Q 0.02fF
C1361 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<26> 0.16fF
C1362 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<14> 0.22fF
C1363 BU_3VX2_16|Q BU_3VX2_9|Q 4.88fF
C1364 BU_3VX2_35|Q BU_3VX2_8|Q 2.81fF
C1365 BU_3VX2_30|Q BU_3VX2_9|Q 2.55fF
C1366 BU_3VX2_69|Q BU_3VX2_22|Q 36.14fF
C1367 BU_3VX2_68|Q BU_3VX2_17|Q 1.99fF
C1368 BU_3VX2_65|Q BU_3VX2_67|Q 13.07fF
C1369 BU_3VX2_18|Q BU_3VX2_7|Q 4.45fF
C1370 BU_3VX2_5|Q BU_3VX2_10|Q 8.05fF
C1371 BU_3VX2_73|Q BU_3VX2_54|Q 0.01fF
C1372 BU_3VX2_42|Q BU_3VX2_50|Q 36.90fF
C1373 BU_3VX2_42|A BU_3VX2_43|Q 0.03fF
C1374 raven_padframe_0|FILLER20F_6|GNDR raven_padframe_0|FILLER20F_6|GNDO 0.81fF
C1375 BU_3VX2_22|A BU_3VX2_26|A 5.71fF
C1376 BU_3VX2_65|A BU_3VX2_64|A 24.61fF
C1377 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<3> 4.09fF
C1378 LS_3VX2_13|A raven_soc_0|ser_rx 0.01fF
C1379 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<9> 0.01fF
C1380 raven_soc_0|flash_io0_do BU_3VX2_33|Q 0.01fF
C1381 AMUX4_3V_1|SEL[1] BU_3VX2_53|Q 36.87fF
C1382 raven_soc_0|gpio_pulldown<7> vdd 0.21fF
C1383 raven_soc_0|ram_wdata<19> apllc03_1v8_0|CLK 0.01fF
C1384 raven_soc_0|irq_pin BU_3VX2_60|Q 0.01fF
C1385 LS_3VX2_21|A LS_3VX2_20|A 58.30fF
C1386 BU_3VX2_22|A BU_3VX2_11|A 1.33fF
C1387 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<12> 0.01fF
C1388 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<15> 0.01fF
C1389 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<7> 0.01fF
C1390 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<9> 4.54fF
C1391 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<6> 2.64fF
C1392 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<11> 0.01fF
C1393 VDD raven_padframe_0|CORNERESDF_2|VDDR 0.71fF
C1394 raven_padframe_0|FILLER20F_8|VDDR raven_padframe_0|FILLER20F_8|GNDR 0.68fF
C1395 LS_3VX2_7|A BU_3VX2_53|Q 9.46fF
C1396 BU_3VX2_31|A VDD3V3 6.11fF
C1397 BU_3VX2_12|A vdd 0.06fF
C1398 BU_3VX2_0|Q raven_soc_0|ram_wdata<18> 0.02fF
C1399 VDD raven_padframe_0|FILLER02F_1|GNDR 0.20fF
C1400 raven_padframe_0|APR00DF_0|VDDR raven_padframe_0|APR00DF_0|GNDR 0.68fF
C1401 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<31> 3.43fF
C1402 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<15> 2.09fF
C1403 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<27> 37.48fF
C1404 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<16> 8.60fF
C1405 raven_soc_0|ram_rdata<30> raven_soc_0|ram_addr<0> 32.52fF
C1406 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<1> 1.89fF
C1407 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<17> 0.01fF
C1408 raven_soc_0|flash_io1_di raven_soc_0|flash_clk 14.83fF
C1409 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<13> 0.01fF
C1410 BU_3VX2_46|A BU_3VX2_44|Q 0.03fF
C1411 raven_padframe_0|GNDORPADF_0|VDDR raven_padframe_0|GNDORPADF_0|GNDOR 0.81fF
C1412 markings_0|date_0|_alphabet_8_0|m2_9_235# markings_0|date_0|_alphabet_0_0|m2_0_208# 0.12fF
C1413 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<15> 0.61fF
C1414 BU_3VX2_9|A raven_soc_0|flash_io1_di 0.01fF
C1415 BU_3VX2_4|A raven_soc_0|flash_io3_oeb 0.01fF
C1416 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<3> 5.11fF
C1417 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<13> 0.01fF
C1418 BU_3VX2_14|A BU_3VX2_12|Q 0.03fF
C1419 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<7> 0.01fF
C1420 raven_soc_0|gpio_in<4> raven_soc_0|ext_clk 0.01fF
C1421 LS_3VX2_4|A BU_3VX2_59|Q 15.66fF
C1422 raven_soc_0|gpio_pullup<11> BU_3VX2_26|Q 0.01fF
C1423 raven_soc_0|gpio_pullup<10> BU_3VX2_25|Q 0.01fF
C1424 raven_soc_0|gpio_pullup<3> apllc03_1v8_0|CLK 0.01fF
C1425 raven_soc_0|gpio_outenb<0> apllc03_1v8_0|B_CP 0.01fF
C1426 raven_soc_0|gpio_pullup<9> BU_3VX2_24|Q 0.01fF
C1427 BU_3VX2_2|A BU_3VX2_4|A 5.65fF
C1428 LS_3VX2_5|Q LS_3VX2_4|Q 2.20fF
C1429 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<8> 0.01fF
C1430 LS_3VX2_3|A raven_soc_0|gpio_outenb<0> 0.01fF
C1431 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<4> 0.01fF
C1432 BU_3VX2_72|A BU_3VX2_29|Q 0.01fF
C1433 BU_3VX2_14|A raven_soc_0|flash_io0_do 0.01fF
C1434 BU_3VX2_63|Q raven_soc_0|flash_io0_di 17.97fF
C1435 LS_3VX2_6|A BU_3VX2_60|Q 0.01fF
C1436 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<9> 4.86fF
C1437 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<13> 0.02fF
C1438 BU_3VX2_40|Q raven_soc_0|gpio_in<6> 0.01fF
C1439 raven_soc_0|ext_clk raven_soc_0|gpio_in<7> 0.01fF
C1440 BU_3VX2_53|A BU_3VX2_60|A 0.41fF
C1441 BU_3VX2_56|A BU_3VX2_57|A 9.03fF
C1442 BU_3VX2_55|A BU_3VX2_58|A 1.50fF
C1443 BU_3VX2_52|A BU_3VX2_61|A 0.25fF
C1444 BU_3VX2_54|A BU_3VX2_59|A 0.71fF
C1445 VDD3V3 LS_3VX2_16|Q 0.44fF
C1446 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<1> 114.65fF
C1447 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<1> 13.27fF
C1448 BU_3VX2_21|A BU_3VX2_26|A 4.37fF
C1449 BU_3VX2_66|A BU_3VX2_65|A 24.75fF
C1450 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<1> 0.01fF
C1451 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<9> 0.01fF
C1452 raven_soc_0|gpio_outenb<2> BU_3VX2_0|Q 0.01fF
C1453 raven_soc_0|gpio_out<10> BU_3VX2_40|Q 0.31fF
C1454 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<11> 0.02fF
C1455 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<9> 1.53fF
C1456 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<8> 2.15fF
C1457 raven_soc_0|gpio_out<8> VDD3V3 0.07fF
C1458 BU_3VX2_21|Q BU_3VX2_23|Q 26.43fF
C1459 BU_3VX2_6|Q BU_3VX2_27|Q 1.08fF
C1460 BU_3VX2_2|Q BU_3VX2_28|Q 21.30fF
C1461 BU_3VX2_13|Q apllc03_1v8_0|CLK 0.01fF
C1462 BU_3VX2_8|Q BU_3VX2_23|Q 2.73fF
C1463 BU_3VX2_17|Q BU_3VX2_24|Q 5.93fF
C1464 BU_3VX2_10|Q BU_3VX2_28|Q 6.66fF
C1465 BU_3VX2_22|Q BU_3VX2_29|Q 4.87fF
C1466 BU_3VX2_7|Q BU_3VX2_27|Q 0.27fF
C1467 BU_3VX2_0|A BU_3VX2_67|A 0.64fF
C1468 BU_3VX2_21|A BU_3VX2_11|A 1.49fF
C1469 LOGIC1_3V_0|Q LOGIC0_3V_2|Q 0.32fF
C1470 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_outenb<2> 7.67fF
C1471 LS_3VX2_8|A AMUX2_3V_0|SEL 32.27fF
C1472 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<10> 0.01fF
C1473 BU_3VX2_10|A BU_3VX2_10|Q 0.08fF
C1474 LS_3VX2_14|A BU_3VX2_73|Q 24.82fF
C1475 LS_3VX2_13|Q VDD3V3 0.16fF
C1476 BU_3VX2_0|Q BU_3VX2_64|Q 0.01fF
C1477 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<18> 0.83fF
C1478 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<24> 52.88fF
C1479 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<21> 0.84fF
C1480 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<14> 4.47fF
C1481 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_outenb<9> 5.00fF
C1482 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pullup<13> 0.02fF
C1483 raven_soc_0|ram_rdata<23> vdd 0.71fF
C1484 raven_soc_0|flash_io2_di BU_3VX2_27|Q 0.01fF
C1485 raven_soc_0|flash_clk BU_3VX2_28|Q 15.69fF
C1486 BU_3VX2_46|A vdd 0.06fF
C1487 LS_3VX2_18|Q VDD3V3 0.57fF
C1488 BU_3VX2_10|A raven_soc_0|flash_clk 0.01fF
C1489 raven_spi_0|SDI raven_soc_0|gpio_out<15> 4.45fF
C1490 BU_3VX2_22|A VDD3V3 0.46fF
C1491 IN_3VX2_1|A raven_soc_0|gpio_in<15> 0.01fF
C1492 raven_soc_0|gpio_in<3> BU_3VX2_40|Q 0.01fF
C1493 raven_padframe_0|ICF_1|VDDR raven_padframe_0|ICF_1|VDDO 0.06fF
C1494 IN_3VX2_1|A BU_3VX2_43|Q 13.04fF
C1495 BU_3VX2_28|A raven_soc_0|flash_io1_di 0.01fF
C1496 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<9> 1.21fF
C1497 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<12> 11.27fF
C1498 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<8> 0.28fF
C1499 LS_3VX2_3|A raven_soc_0|flash_io0_do 0.01fF
C1500 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<13> 16.64fF
C1501 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<15> 0.02fF
C1502 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<10> 5.95fF
C1503 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<7> 0.01fF
C1504 raven_soc_0|gpio_out<9> BU_3VX2_40|Q 0.01fF
C1505 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<6> 3.95fF
C1506 raven_soc_0|gpio_out<7> raven_soc_0|ext_clk 0.01fF
C1507 raven_soc_0|gpio_out<6> VDD3V3 0.27fF
C1508 raven_padframe_0|BBCUD4F_3|VDDR raven_padframe_0|BBCUD4F_3|VDDO 0.06fF
C1509 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<20> 4.27fF
C1510 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<0> 2.19fF
C1511 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<19> 0.02fF
C1512 LS_3VX2_21|A BU_3VX2_47|Q 13.38fF
C1513 BU_3VX2_10|A BU_3VX2_9|A 31.49fF
C1514 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<3> 3.25fF
C1515 LS_3VX2_12|Q LS_3VX2_7|Q 15.11fF
C1516 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<3> 0.01fF
C1517 BU_3VX2_0|A raven_soc_0|flash_clk 0.01fF
C1518 BU_3VX2_5|A raven_soc_0|flash_io0_di 0.04fF
C1519 LS_3VX2_8|A BU_3VX2_61|Q 0.01fF
C1520 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<5> 0.01fF
C1521 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<13> 14.14fF
C1522 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<8> 2.11fF
C1523 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<10> 0.23fF
C1524 raven_soc_0|ram_wenb raven_soc_0|ram_addr<8> 0.01fF
C1525 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pulldown<6> 0.03fF
C1526 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pullup<13> 6.65fF
C1527 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<14> 0.02fF
C1528 VDD raven_padframe_0|BBCUD4F_1|VDDR 0.71fF
C1529 raven_soc_0|gpio_pulldown<8> BU_3VX2_26|Q 0.01fF
C1530 raven_soc_0|gpio_pulldown<11> BU_3VX2_27|Q 0.01fF
C1531 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<3> 0.08fF
C1532 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<15> 7.82fF
C1533 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<12> 0.02fF
C1534 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<14> 3.42fF
C1535 BU_3VX2_73|Q BU_3VX2_56|Q 0.01fF
C1536 BU_3VX2_64|Q BU_3VX2_30|Q 16.84fF
C1537 BU_3VX2_31|Q BU_3VX2_69|Q 1.53fF
C1538 AMUX4_3V_4|SEL[1] BU_3VX2_7|Q 0.01fF
C1539 LS_3VX2_27|Q BU_3VX2_42|Q 0.23fF
C1540 BU_3VX2_42|Q BU_3VX2_48|Q 23.22fF
C1541 raven_padframe_0|FILLER20F_1|GNDR raven_padframe_0|FILLER20F_1|GNDO 0.81fF
C1542 BU_3VX2_23|A BU_3VX2_18|A 4.50fF
C1543 BU_3VX2_9|A BU_3VX2_0|A 0.01fF
C1544 LS_3VX2_11|Q LS_3VX2_7|A 0.54fF
C1545 analog_out adc_low 0.38fF
C1546 raven_padframe_0|BBCUD4F_7|GNDR raven_padframe_0|BBCUD4F_7|GNDO 0.81fF
C1547 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<5> 0.80fF
C1548 LS_3VX2_4|A AMUX2_3V_0|SEL 8.15fF
C1549 raven_soc_0|gpio_pulldown<14> LS_3VX2_3|A 0.01fF
C1550 raven_padframe_0|CORNERESDF_1|VDDR raven_padframe_0|CORNERESDF_1|GNDR 0.68fF
C1551 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<0> 12.02fF
C1552 raven_soc_0|flash_io1_di BU_3VX2_33|Q 0.01fF
C1553 raven_soc_0|ram_wdata<21> vdd 0.98fF
C1554 raven_soc_0|ram_wdata<30> apllc03_1v8_0|CLK 0.01fF
C1555 raven_soc_0|irq_pin BU_3VX2_62|Q 0.01fF
C1556 LS_3VX2_27|A LS_3VX2_20|A 35.35fF
C1557 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<12> 0.97fF
C1558 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<5> 0.04fF
C1559 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<12> 0.01fF
C1560 IN_3VX2_1|A raven_soc_0|gpio_out<13> 0.01fF
C1561 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<7> 0.01fF
C1562 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<6> 25.68fF
C1563 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<9> 3.31fF
C1564 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<5> 0.02fF
C1565 raven_soc_0|gpio_out<2> BU_3VX2_63|Q 0.01fF
C1566 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<11> 0.01fF
C1567 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<7> 0.01fF
C1568 BU_3VX2_33|A raven_soc_0|gpio_pulldown<15> 2.26fF
C1569 BU_3VX2_6|A BU_3VX2_6|Q 0.08fF
C1570 BU_3VX2_6|A BU_3VX2_7|Q 0.03fF
C1571 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<5> 0.07fF
C1572 LS_3VX2_24|A BU_3VX2_42|Q 13.29fF
C1573 raven_soc_0|gpio_pulldown<2> VDD3V3 3.51fF
C1574 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<30> 3.10fF
C1575 raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<4> 14.36fF
C1576 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<31> 63.67fF
C1577 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<20> 0.01fF
C1578 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<24> 0.01fF
C1579 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io2_di 25.29fF
C1580 BU_3VX2_36|Q BU_3VX2_67|Q 4.21fF
C1581 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<31> 5.62fF
C1582 BU_3VX2_21|Q BU_3VX2_4|Q 12.13fF
C1583 BU_3VX2_4|Q BU_3VX2_8|Q 13.38fF
C1584 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<26> 61.37fF
C1585 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<17> 4.15fF
C1586 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<13> 5.73fF
C1587 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<1> 1.45fF
C1588 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io0_oeb 92.96fF
C1589 raven_soc_0|flash_io1_do raven_soc_0|flash_io0_do 375.23fF
C1590 BU_3VX2_38|Q BU_3VX2_36|Q 0.02fF
C1591 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<17> 0.05fF
C1592 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<21> 0.38fF
C1593 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<25> 0.01fF
C1594 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<22> 0.01fF
C1595 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<27> 2.59fF
C1596 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<19> 2.88fF
C1597 BU_3VX2_59|Q vdd 2.31fF
C1598 raven_padframe_0|FILLER20F_5|GNDR raven_padframe_0|FILLER20F_5|GNDO 0.81fF
C1599 BU_3VX2_6|A raven_soc_0|flash_io2_di 0.03fF
C1600 BU_3VX2_2|A raven_soc_0|flash_io0_oeb 0.01fF
C1601 BU_3VX2_21|A VDD3V3 0.33fF
C1602 IN_3VX2_1|Q BU_3VX2_53|Q 0.01fF
C1603 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<6> 0.45fF
C1604 BU_3VX2_28|A BU_3VX2_28|Q 0.08fF
C1605 raven_padframe_0|BBCUD4F_13|VDDR raven_padframe_0|BBCUD4F_13|VDDO 0.06fF
C1606 IN_3VX2_1|A BU_3VX2_50|Q 0.01fF
C1607 LS_3VX2_4|A BU_3VX2_61|Q 7.14fF
C1608 raven_soc_0|gpio_pullup<4> vdd 0.40fF
C1609 raven_soc_0|gpio_pulldown<5> apllc03_1v8_0|CLK 0.03fF
C1610 raven_soc_0|gpio_pulldown<9> BU_3VX2_24|Q 0.01fF
C1611 BU_3VX2_71|Q raven_soc_0|flash_io1_oeb 0.40fF
C1612 BU_3VX2_10|A BU_3VX2_28|A 0.01fF
C1613 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<7> 0.01fF
C1614 LS_3VX2_3|A raven_soc_0|gpio_pulldown<10> 0.01fF
C1615 BU_3VX2_35|A raven_soc_0|flash_io3_do 0.09fF
C1616 VDD raven_padframe_0|BBC4F_2|GNDO 0.07fF
C1617 VDD raven_padframe_0|FILLER10F_1|GNDR 0.16fF
C1618 BU_3VX2_67|A vdd 0.22fF
C1619 VDD raven_padframe_0|BBCUD4F_14|GNDO 0.07fF
C1620 BU_3VX2_14|A raven_soc_0|flash_io1_di 0.01fF
C1621 AMUX2_3V_0|SEL comp_inp 1.13fF
C1622 LS_3VX2_13|A AMUX4_3V_1|SEL[0] 8.11fF
C1623 LS_3VX2_6|A BU_3VX2_62|Q 0.01fF
C1624 BU_3VX2_40|Q raven_soc_0|ext_clk 100.17fF
C1625 LS_3VX2_27|Q BU_3VX2_42|A 2.81fF
C1626 VDD3V3 BU_3VX2_53|A 0.05fF
C1627 raven_padframe_0|POWERCUTVDD3FC_0|GNDR raven_padframe_0|POWERCUTVDD3FC_0|GNDO 0.77fF
C1628 BU_3VX2_0|A BU_3VX2_28|A 0.01fF
C1629 BU_3VX2_18|A IN_3VX2_1|A 1.77fF
C1630 raven_padframe_0|BBCUD4F_3|VDDO raven_padframe_0|BBCUD4F_3|GNDO 2.28fF
C1631 LS_3VX2_5|A LS_3VX2_6|A 55.76fF
C1632 BU_3VX2_31|A raven_soc_0|gpio_pullup<8> 0.01fF
C1633 raven_padframe_0|GNDORPADF_1|VDDR raven_padframe_0|GNDORPADF_1|VDDO 0.06fF
C1634 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<4> 0.16fF
C1635 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_outenb<6> 0.25fF
C1636 markings_0|product_name_0|_alphabet_V_0|m2_0_560# markings_0|product_name_0|_alphabet_R_0|m2_0_0# 0.09fF
C1637 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<13> 0.02fF
C1638 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<14> 15.84fF
C1639 raven_soc_0|gpio_pulldown<6> VDD3V3 0.07fF
C1640 BU_3VX2_35|Q BU_3VX2_27|Q 0.01fF
C1641 BU_3VX2_19|Q BU_3VX2_23|Q 9.57fF
C1642 BU_3VX2_18|Q BU_3VX2_23|Q 12.24fF
C1643 BU_3VX2_9|Q BU_3VX2_26|Q 7.56fF
C1644 BU_3VX2_2|Q vdd 1.60fF
C1645 BU_3VX2_10|Q vdd 1.03fF
C1646 BU_3VX2_31|Q BU_3VX2_29|Q 22.87fF
C1647 BU_3VX2_7|Q BU_3VX2_25|Q 0.22fF
C1648 BU_3VX2_6|Q BU_3VX2_25|Q 0.27fF
C1649 BU_3VX2_69|Q apllc03_1v8_0|CLK 0.01fF
C1650 raven_soc_0|irq_pin BU_3VX2_45|Q 15.54fF
C1651 BU_3VX2_15|Q BU_3VX2_26|Q 3.21fF
C1652 BU_3VX2_23|A BU_3VX2_71|A 0.01fF
C1653 raven_padframe_0|ICFC_2|VDDR LOGIC0_3V_4|Q 0.01fF
C1654 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<3> 0.01fF
C1655 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<10> 0.01fF
C1656 BU_3VX2_70|A BU_3VX2_69|Q 0.16fF
C1657 raven_soc_0|ram_rdata<13> raven_soc_0|ram_rdata<17> 15.74fF
C1658 raven_soc_0|ram_wdata<27> raven_soc_0|ram_rdata<16> 0.38fF
C1659 raven_soc_0|ram_rdata<1> raven_soc_0|ram_addr<0> 0.02fF
C1660 raven_soc_0|ram_wdata<31> raven_soc_0|ram_rdata<15> 0.01fF
C1661 raven_soc_0|flash_clk vdd 2.84fF
C1662 raven_soc_0|flash_io3_oeb BU_3VX2_29|Q 0.01fF
C1663 raven_soc_0|flash_io0_di BU_3VX2_24|Q 0.01fF
C1664 raven_soc_0|flash_io0_oeb apllc03_1v8_0|CLK 0.01fF
C1665 raven_soc_0|flash_io2_di BU_3VX2_25|Q 0.01fF
C1666 raven_padframe_0|FILLER01F_1|VDDR raven_padframe_0|FILLER01F_1|GNDO 0.13fF
C1667 raven_padframe_0|BBC4F_3|VDDO raven_padframe_0|BBC4F_3|GNDO 2.28fF
C1668 raven_padframe_0|axtoc02_3v3_0|m4_0_28769# raven_padframe_0|axtoc02_3v3_0|GNDO 0.07fF
C1669 raven_padframe_0|axtoc02_3v3_0|m4_55000_30653# raven_padframe_0|axtoc02_3v3_0|VDDR 0.15fF
C1670 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<5> 0.01fF
C1671 BU_3VX2_3|A raven_soc_0|ext_clk 0.01fF
C1672 BU_3VX2_9|A vdd 0.11fF
C1673 BU_3VX2_15|A raven_soc_0|ext_clk 0.01fF
C1674 VDD raven_padframe_0|FILLER20F_8|GNDR 0.16fF
C1675 IN_3VX2_1|A raven_soc_0|gpio_in<14> 0.01fF
C1676 adc_high raven_soc_0|ser_tx 0.13fF
C1677 VDD raven_padframe_0|BBCUD4F_5|GNDO 0.07fF
C1678 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pullup<5> 1.49fF
C1679 LS_3VX2_3|A raven_soc_0|flash_io1_di 0.12fF
C1680 BU_3VX2_0|Q raven_soc_0|flash_io3_do 0.20fF
C1681 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<7> 0.01fF
C1682 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<8> 0.01fF
C1683 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<13> 39.36fF
C1684 raven_soc_0|gpio_outenb<10> BU_3VX2_40|Q 0.01fF
C1685 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<15> 0.02fF
C1686 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<12> 0.01fF
C1687 raven_soc_0|gpio_outenb<11> VDD3V3 0.07fF
C1688 raven_soc_0|gpio_outenb<7> raven_soc_0|ext_clk 0.01fF
C1689 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<6> 0.01fF
C1690 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<19> 0.20fF
C1691 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<23> 150.13fF
C1692 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<0> 1.52fF
C1693 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<20> 0.01fF
C1694 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<11> 0.01fF
C1695 LS_3VX2_27|A BU_3VX2_47|Q 12.31fF
C1696 LS_3VX2_12|Q LS_3VX2_4|Q 0.52fF
C1697 BU_3VX2_40|A raven_soc_0|flash_clk 0.01fF
C1698 VDD raven_padframe_0|BT4F_0|GNDR 0.16fF
C1699 LS_3VX2_8|A LS_3VX2_15|A 0.02fF
C1700 BU_3VX2_13|A raven_soc_0|flash_io0_di 0.01fF
C1701 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<13> 12.82fF
C1702 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_outenb<9> 0.13fF
C1703 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<3> 0.08fF
C1704 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<27> 0.16fF
C1705 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<5> 0.01fF
C1706 BU_3VX2_27|A raven_soc_0|flash_io2_di 0.01fF
C1707 BU_3VX2_0|Q raven_soc_0|gpio_out<14> 0.01fF
C1708 BU_3VX2_33|A raven_soc_0|flash_io3_di 0.22fF
C1709 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<8> 11.28fF
C1710 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pulldown<6> 10.94fF
C1711 raven_soc_0|gpio_pulldown<13> BU_3VX2_71|Q 0.01fF
C1712 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pulldown<7> 0.02fF
C1713 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<8> 0.88fF
C1714 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<10> 111.23fF
C1715 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<13> 2.51fF
C1716 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<14> 2.89fF
C1717 AMUX2_3V_0|SEL vdd 3.03fF
C1718 raven_soc_0|gpio_pulldown<11> BU_3VX2_25|Q 0.01fF
C1719 BU_3VX2_63|Q BU_3VX2_24|Q 0.01fF
C1720 LS_3VX2_13|A LS_3VX2_17|A 0.01fF
C1721 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<11> 6.15fF
C1722 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<1> 2.78fF
C1723 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<0> 1.68fF
C1724 LS_3VX2_20|Q LS_3VX2_20|A 0.06fF
C1725 BU_3VX2_7|A BU_3VX2_17|A 1.14fF
C1726 BU_3VX2_9|A BU_3VX2_40|A 0.51fF
C1727 BU_3VX2_19|A BU_3VX2_31|A 1.73fF
C1728 BU_3VX2_10|A BU_3VX2_14|A 3.38fF
C1729 raven_padframe_0|APR00DF_3|VDDR raven_padframe_0|APR00DF_3|GNDR 0.68fF
C1730 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<14> 15.54fF
C1731 raven_padframe_0|BT4F_0|VDDR raven_padframe_0|BT4F_0|GNDO 0.13fF
C1732 raven_soc_0|gpio_pullup<1> BU_3VX2_71|Q 0.07fF
C1733 LOGIC0_3V_4|Q raven_padframe_0|ICF_2|PO 0.04fF
C1734 raven_soc_0|ram_rdata<3> vdd 0.28fF
C1735 LS_3VX2_19|A VDD3V3 0.74fF
C1736 raven_soc_0|ram_wdata<14> vdd 0.72fF
C1737 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<12> 0.01fF
C1738 BU_3VX2_8|A BU_3VX2_35|A 0.72fF
C1739 BU_3VX2_25|A BU_3VX2_18|A 3.12fF
C1740 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<7> 0.01fF
C1741 BU_3VX2_71|A IN_3VX2_1|A 0.01fF
C1742 BU_3VX2_0|A BU_3VX2_14|A 0.01fF
C1743 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<15> 0.01fF
C1744 IN_3VX2_1|A raven_soc_0|gpio_outenb<15> 0.01fF
C1745 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<0> 149.98fF
C1746 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<9> 0.01fF
C1747 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<11> 0.56fF
C1748 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<12> 0.34fF
C1749 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<10> 1.02fF
C1750 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<6> 0.01fF
C1751 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<12> 0.02fF
C1752 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<9> 14.98fF
C1753 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<7> 0.01fF
C1754 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<5> 0.01fF
C1755 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<30> 180.40fF
C1756 raven_soc_0|flash_io1_do raven_soc_0|flash_io1_di 82.07fF
C1757 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<24> 28.31fF
C1758 raven_soc_0|flash_io2_do raven_soc_0|flash_io3_oeb 81.05fF
C1759 BU_3VX2_19|Q BU_3VX2_4|Q 2.19fF
C1760 BU_3VX2_15|Q BU_3VX2_11|Q 13.85fF
C1761 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<27> 0.08fF
C1762 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<10> 0.05fF
C1763 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<25> 15.68fF
C1764 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<15> 3.85fF
C1765 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<2> 6.76fF
C1766 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<14> 0.09fF
C1767 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<26> 0.02fF
C1768 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<19> 0.02fF
C1769 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<8> 1.48fF
C1770 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<6> 8.78fF
C1771 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<8> 0.01fF
C1772 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<4> 5.76fF
C1773 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<22> 0.21fF
C1774 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<25> 0.11fF
C1775 raven_soc_0|flash_io3_do raven_soc_0|flash_io3_di 322.52fF
C1776 BU_3VX2_2|Q BU_3VX2_70|Q 0.01fF
C1777 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<29> 3.16fF
C1778 AMUX4_3V_3|SEL[1] LS_3VX2_18|A 0.85fF
C1779 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<2> 0.01fF
C1780 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<21> 0.01fF
C1781 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<17> 0.01fF
C1782 AMUX4_3V_4|SEL[0] BU_3VX2_33|Q 31.10fF
C1783 BU_3VX2_36|Q BU_3VX2_65|Q 7.96fF
C1784 BU_3VX2_4|Q BU_3VX2_18|Q 0.87fF
C1785 BU_3VX2_3|Q BU_3VX2_8|Q 21.49fF
C1786 BU_3VX2_70|Q BU_3VX2_10|Q 2.64fF
C1787 BU_3VX2_11|Q BU_3VX2_9|Q 23.99fF
C1788 BU_3VX2_23|Q BU_3VX2_27|Q 59.29fF
C1789 BU_3VX2_61|Q vdd 2.53fF
C1790 BU_3VX2_28|Q apllc03_1v8_0|B_CP 0.61fF
C1791 apllc03_1v8_0|CLK BU_3VX2_29|Q 10.20fF
C1792 raven_soc_0|gpio_in<11> raven_padframe_0|BBCUD4F_11|PO 0.04fF
C1793 raven_padframe_0|ICFC_0|VDDR LOGIC0_3V_4|Q 0.01fF
C1794 raven_padframe_0|FILLER50F_1|VDDO raven_padframe_0|FILLER50F_1|GNDO 2.28fF
C1795 raven_padframe_0|BBCUD4F_12|GNDR raven_padframe_0|BBCUD4F_12|VDDO 0.09fF
C1796 BU_3VX2_2|A raven_soc_0|flash_io2_do 0.01fF
C1797 BU_3VX2_38|A raven_soc_0|flash_io2_oeb 0.01fF
C1798 adc_low VDD3V3 27.57fF
C1799 IN_3VX2_1|A BU_3VX2_48|Q 6.20fF
C1800 BU_3VX2_28|A vdd 0.06fF
C1801 VDD raven_padframe_0|FILLER20F_4|GNDR 0.16fF
C1802 LS_3VX2_4|A LS_3VX2_15|A 6.56fF
C1803 LS_3VX2_3|A BU_3VX2_28|Q 0.01fF
C1804 raven_soc_0|ser_rx LS_3VX2_17|A 10.43fF
C1805 raven_soc_0|gpio_in<5> raven_soc_0|flash_io0_di 0.15fF
C1806 BU_3VX2_6|A BU_3VX2_38|A 1.28fF
C1807 BU_3VX2_7|A BU_3VX2_12|A 2.39fF
C1808 BU_3VX2_22|A BU_3VX2_21|Q 0.16fF
C1809 raven_soc_0|gpio_pulldown<12> LS_3VX2_3|A 0.01fF
C1810 LS_3VX2_8|A AMUX4_3V_1|SEL[1] 9.22fF
C1811 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<12> 0.01fF
C1812 BU_3VX2_63|Q raven_soc_0|gpio_out<15> 0.06fF
C1813 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<10> 0.01fF
C1814 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<8> 74.43fF
C1815 raven_soc_0|gpio_outenb<2> BU_3VX2_26|Q 0.01fF
C1816 raven_soc_0|gpio_out<2> BU_3VX2_24|Q 0.01fF
C1817 LS_3VX2_8|A LS_3VX2_7|A 52.88fF
C1818 BU_3VX2_40|A BU_3VX2_28|A 0.02fF
C1819 raven_soc_0|gpio_pulldown<1> BU_3VX2_0|Q 0.16fF
C1820 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<13> 0.01fF
C1821 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<8> 0.48fF
C1822 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<12> 3.50fF
C1823 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<13> 0.02fF
C1824 BU_3VX2_63|Q raven_soc_0|gpio_in<5> 0.01fF
C1825 raven_soc_0|flash_csb raven_soc_0|flash_io0_do 41.01fF
C1826 BU_3VX2_24|A BU_3VX2_23|A 63.03fF
C1827 LOGIC0_3V_1|Q LOGIC1_3V_1|Q 0.51fF
C1828 raven_soc_0|flash_io3_do raven_soc_0|irq_pin 0.01fF
C1829 raven_soc_0|irq_pin AMUX4_3V_4|AIN3 42.60fF
C1830 BU_3VX2_64|Q BU_3VX2_26|Q 3.58fF
C1831 BU_3VX2_68|Q BU_3VX2_24|Q 1.37fF
C1832 BU_3VX2_33|Q vdd 1.49fF
C1833 BU_3VX2_35|Q BU_3VX2_25|Q 0.01fF
C1834 BU_3VX2_22|A BU_3VX2_19|A 7.27fF
C1835 VDD raven_padframe_0|BBCUD4F_3|VDDR 0.71fF
C1836 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<4> 1.68fF
C1837 BU_3VX2_5|A BU_3VX2_13|A 1.34fF
C1838 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<0> 17.33fF
C1839 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<1> 3.26fF
C1840 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<4> 5.44fF
C1841 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<16> 0.02fF
C1842 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<0> 8.29fF
C1843 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<17> 0.01fF
C1844 raven_soc_0|ram_wdata<19> raven_soc_0|ram_rdata<15> 2.10fF
C1845 raven_soc_0|ram_wdata<29> raven_soc_0|ram_rdata<1> 5.89fF
C1846 raven_soc_0|ram_wdata<26> raven_soc_0|ram_rdata<16> 0.27fF
C1847 raven_soc_0|ram_wdata<22> raven_soc_0|ram_rdata<13> 0.46fF
C1848 BU_3VX2_45|A LS_3VX2_20|Q 0.49fF
C1849 BU_3VX2_41|A BU_3VX2_42|A 0.21fF
C1850 BU_3VX2_46|A LS_3VX2_21|Q 0.25fF
C1851 BU_3VX2_60|A BU_3VX2_60|Q 0.10fF
C1852 BU_3VX2_48|A BU_3VX2_49|Q 0.03fF
C1853 BU_3VX2_51|A BU_3VX2_50|Q 0.15fF
C1854 raven_soc_0|flash_io2_do apllc03_1v8_0|CLK 11.38fF
C1855 raven_soc_0|flash_io2_oeb BU_3VX2_23|Q 0.01fF
C1856 BU_3VX2_62|A BU_3VX2_61|Q 0.03fF
C1857 raven_soc_0|flash_io1_do BU_3VX2_28|Q 0.01fF
C1858 BU_3VX2_25|A BU_3VX2_71|A 0.01fF
C1859 raven_padframe_0|FILLER01F_0|VDDR raven_padframe_0|FILLER01F_0|VDDO 0.06fF
C1860 raven_padframe_0|BBCUD4F_3|VDDR LOGIC0_3V_4|Q 0.01fF
C1861 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<15> 0.01fF
C1862 raven_padframe_0|aregc01_3v3_1|m4_92500_29057# raven_padframe_0|aregc01_3v3_1|VDDO 0.04fF
C1863 raven_padframe_0|aregc01_3v3_1|m4_92500_29333# raven_padframe_0|aregc01_3v3_1|GNDO 0.12fF
C1864 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<14> 0.01fF
C1865 raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# raven_padframe_0|axtoc02_3v3_0|m4_55000_28769# 0.02fF
C1866 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<12> 0.01fF
C1867 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<5> 0.01fF
C1868 BU_3VX2_10|A raven_soc_0|flash_io1_do 0.03fF
C1869 BU_3VX2_63|A raven_soc_0|flash_io3_do 0.01fF
C1870 LS_3VX2_10|A BU_3VX2_54|Q 10.83fF
C1871 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<6> 0.01fF
C1872 LS_3VX2_4|A AMUX4_3V_1|SEL[1] 158.61fF
C1873 AMUX2_3V_0|AOUT VDD3V3 2.94fF
C1874 raven_soc_0|gpio_pullup<10> BU_3VX2_40|Q 0.37fF
C1875 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<5> 2.86fF
C1876 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<15> 0.02fF
C1877 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<10> 123.60fF
C1878 raven_soc_0|gpio_pullup<9> raven_soc_0|ext_clk 0.01fF
C1879 raven_soc_0|gpio_pullup<11> VDD3V3 0.07fF
C1880 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<0> 0.01fF
C1881 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<20> 0.22fF
C1882 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<11> 4.23fF
C1883 raven_soc_0|gpio_outenb<8> BU_3VX2_29|Q 0.01fF
C1884 BU_3VX2_4|Q BU_3VX2_27|Q 4.57fF
C1885 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<4> 0.05fF
C1886 LS_3VX2_7|A LS_3VX2_4|A 14.74fF
C1887 BU_3VX2_21|A BU_3VX2_21|Q 0.08fF
C1888 BU_3VX2_8|A raven_soc_0|flash_io3_di 0.01fF
C1889 BU_3VX2_20|A raven_soc_0|flash_io0_do 0.01fF
C1890 BU_3VX2_0|A raven_soc_0|flash_io1_do 5.74fF
C1891 LOGIC0_3V_4|Q raven_soc_0|gpio_in<9> 0.08fF
C1892 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<14> 21.71fF
C1893 raven_spi_0|sdo_enb raven_soc_0|flash_io0_oeb 0.45fF
C1894 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<10> 39.40fF
C1895 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<6> 0.74fF
C1896 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<11> 4.31fF
C1897 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<12> 2.83fF
C1898 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pulldown<6> 2.61fF
C1899 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pulldown<7> 0.02fF
C1900 BU_3VX2_14|A vdd 0.06fF
C1901 raven_padframe_0|BBCUD4F_0|VDDR raven_padframe_0|BBCUD4F_0|GNDR 0.68fF
C1902 raven_spi_0|SDO BU_3VX2_33|A 29.71fF
C1903 BU_3VX2_4|A BU_3VX2_18|A 0.01fF
C1904 BU_3VX2_38|A BU_3VX2_27|A 0.01fF
C1905 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<13> 0.62fF
C1906 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<14> 1.29fF
C1907 raven_padframe_0|BBCUD4F_11|VDDR raven_padframe_0|BBCUD4F_11|GNDO 0.13fF
C1908 LS_3VX2_22|A VDD3V3 0.81fF
C1909 raven_soc_0|ram_wdata<11> vdd 0.53fF
C1910 BU_3VX2_24|A IN_3VX2_1|A 6.21fF
C1911 BU_3VX2_56|Q BU_3VX2_43|Q 0.20fF
C1912 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<12> 0.01fF
C1913 BU_3VX2_21|A BU_3VX2_19|A 12.66fF
C1914 BU_3VX2_23|A BU_3VX2_16|A 3.05fF
C1915 BU_3VX2_23|A BU_3VX2_29|A 6.42fF
C1916 LS_3VX2_11|A LS_3VX2_6|A 154.81fF
C1917 raven_soc_0|gpio_out<0> BU_3VX2_0|Q 0.01fF
C1918 LS_3VX2_13|Q LS_3VX2_24|Q 0.01fF
C1919 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<10> 0.01fF
C1920 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<9> 0.01fF
C1921 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<7> 0.09fF
C1922 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<11> 4.46fF
C1923 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<6> 0.16fF
C1924 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<5> 0.02fF
C1925 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<12> 0.02fF
C1926 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<9> 20.84fF
C1927 BU_3VX2_0|Q raven_soc_0|gpio_out<12> 0.01fF
C1928 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<13> 0.02fF
C1929 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<10> 41.69fF
C1930 raven_soc_0|gpio_out<1> apllc03_1v8_0|CLK 0.01fF
C1931 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<6> 14.64fF
C1932 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<4> 4.55fF
C1933 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<7> 0.39fF
C1934 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<18> 9.48fF
C1935 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<6> 0.10fF
C1936 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<5> 0.10fF
C1937 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<8> 3.98fF
C1938 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<31> 0.06fF
C1939 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<22> 4.82fF
C1940 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<20> 21.09fF
C1941 LOGIC0_3V_0|Q LOGIC1_3V_0|Q 0.52fF
C1942 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<3> 0.01fF
C1943 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<2> 2.93fF
C1944 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<12> 0.25fF
C1945 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<26> 0.02fF
C1946 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<25> 19.27fF
C1947 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<14> 0.05fF
C1948 BU_3VX2_19|Q BU_3VX2_3|Q 1.13fF
C1949 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<1> 5.74fF
C1950 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<17> 7.23fF
C1951 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<0> 0.04fF
C1952 BU_3VX2_12|Q BU_3VX2_14|Q 26.44fF
C1953 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<13> 0.53fF
C1954 BU_3VX2_6|Q BU_3VX2_37|Q 9.13fF
C1955 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<15> 7.07fF
C1956 BU_3VX2_3|Q BU_3VX2_18|Q 6.94fF
C1957 BU_3VX2_32|Q BU_3VX2_31|Q 1.03fF
C1958 BU_3VX2_70|Q BU_3VX2_33|Q 0.55fF
C1959 BU_3VX2_37|Q BU_3VX2_7|Q 6.31fF
C1960 raven_soc_0|irq_pin LS_3VX2_21|A 0.01fF
C1961 LS_3VX2_15|A vdd 3.80fF
C1962 BU_3VX2_25|Q BU_3VX2_23|Q 134.71fF
C1963 BU_3VX2_26|Q apllc03_1v8_0|B_VCO 0.98fF
C1964 vdd apllc03_1v8_0|B_CP 3.41fF
C1965 BU_3VX2_23|A BU_3VX2_37|A 0.01fF
C1966 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<0> 29.90fF
C1967 BU_3VX2_67|A BU_3VX2_69|A 8.49fF
C1968 raven_padframe_0|CORNERESDF_0|VDDR raven_padframe_0|CORNERESDF_0|GNDR 0.68fF
C1969 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<11> 0.01fF
C1970 raven_padframe_0|aregc01_3v3_0|GNDR raven_padframe_0|aregc01_3v3_0|GNDO 0.59fF
C1971 raven_padframe_0|BBCUD4F_2|VDDO raven_padframe_0|BBCUD4F_2|GNDO 2.28fF
C1972 raven_spi_0|SDO raven_soc_0|flash_io3_do 0.71fF
C1973 LS_3VX2_14|A BU_3VX2_50|Q 5.59fF
C1974 VDD raven_padframe_0|BBCUD4F_3|GNDO 0.07fF
C1975 BU_3VX2_36|A BU_3VX2_64|Q 0.03fF
C1976 LS_3VX2_3|A vdd 1.09fF
C1977 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<27> 0.01fF
C1978 raven_soc_0|ram_rdata<28> raven_soc_0|ram_addr<0> 14.23fF
C1979 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<17> 14.76fF
C1980 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<31> 0.02fF
C1981 raven_soc_0|ram_wdata<24> apllc03_1v8_0|CLK 0.01fF
C1982 BU_3VX2_22|A BU_3VX2_19|Q 0.02fF
C1983 BU_3VX2_6|A BU_3VX2_4|Q 0.03fF
C1984 VDD raven_padframe_0|BBC4F_3|GNDO 0.07fF
C1985 BU_3VX2_11|A BU_3VX2_9|Q 0.03fF
C1986 BU_3VX2_63|Q raven_soc_0|gpio_in<6> 0.01fF
C1987 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<13> 19.75fF
C1988 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<7> 0.01fF
C1989 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<5> 0.01fF
C1990 BU_3VX2_31|A BU_3VX2_27|Q 32.69fF
C1991 raven_soc_0|gpio_pulldown<8> VDD3V3 0.07fF
C1992 LS_3VX2_13|A BU_3VX2_42|Q 6.98fF
C1993 BU_3VX2_8|A BU_3VX2_63|A 0.02fF
C1994 VDD raven_padframe_0|ICF_2|VDDR 0.71fF
C1995 LS_3VX2_10|A LS_3VX2_14|A 13.26fF
C1996 LS_3VX2_13|Q LS_3VX2_6|Q 1.41fF
C1997 BU_3VX2_40|A LS_3VX2_3|A 1.69fF
C1998 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<0> 17.26fF
C1999 raven_soc_0|gpio_in<2> LS_3VX2_3|A 0.01fF
C2000 raven_soc_0|gpio_in<0> raven_soc_0|flash_io1_di 0.47fF
C2001 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<7> 0.01fF
C2002 raven_soc_0|gpio_in<3> raven_soc_0|flash_io0_di 0.45fF
C2003 BU_3VX2_63|Q raven_soc_0|gpio_out<10> 0.38fF
C2004 raven_soc_0|flash_csb raven_soc_0|flash_io1_di 13.53fF
C2005 LS_3VX2_6|A LS_3VX2_21|A 4.91fF
C2006 BU_3VX2_73|Q AMUX4_3V_4|AIN2 7.19fF
C2007 BU_3VX2_55|Q BU_3VX2_49|Q 0.03fF
C2008 AMUX4_3V_0|SEL[1] BU_3VX2_57|Q 0.69fF
C2009 LS_3VX2_13|Q LS_3VX2_8|Q 17.95fF
C2010 BU_3VX2_23|A LS_3VX2_3|Q 0.01fF
C2011 BU_3VX2_4|A BU_3VX2_71|A 0.01fF
C2012 raven_padframe_0|ICF_2|VDDR LOGIC0_3V_4|Q 0.01fF
C2013 raven_padframe_0|ICFC_0|VDD3 LOGIC0_3V_4|Q 0.05fF
C2014 BU_3VX2_16|A IN_3VX2_1|A 0.01fF
C2015 IN_3VX2_1|A BU_3VX2_29|A 90.07fF
C2016 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<0> 0.01fF
C2017 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<8> 86.63fF
C2018 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<9> 13.38fF
C2019 BU_3VX2_24|A BU_3VX2_25|A 57.33fF
C2020 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<13> 0.61fF
C2021 raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<27> 15.83fF
C2022 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<15> 0.40fF
C2023 raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<17> 0.06fF
C2024 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<16> 0.01fF
C2025 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<22> 0.01fF
C2026 BU_3VX2_66|Q BU_3VX2_1|Q 0.52fF
C2027 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<29> 0.01fF
C2028 raven_soc_0|flash_io1_do vdd 2.36fF
C2029 AMUX4_3V_1|SEL[0] LS_3VX2_17|A 0.05fF
C2030 BU_3VX2_50|A LS_3VX2_20|Q 0.15fF
C2031 BU_3VX2_49|A BU_3VX2_44|A 0.48fF
C2032 BU_3VX2_51|A LS_3VX2_27|Q 0.09fF
C2033 BU_3VX2_60|A BU_3VX2_62|Q 0.03fF
C2034 raven_soc_0|gpio_in<10> BU_3VX2_28|Q 0.01fF
C2035 raven_soc_0|gpio_in<15> BU_3VX2_29|Q 0.01fF
C2036 raven_soc_0|ser_tx BU_3VX2_54|Q 5.08fF
C2037 raven_soc_0|flash_io3_do BU_3VX2_26|Q 0.01fF
C2038 raven_soc_0|gpio_out<15> BU_3VX2_24|Q 0.01fF
C2039 AMUX4_3V_1|SEL[1] vdd 5.43fF
C2040 BU_3VX2_51|A BU_3VX2_48|Q 0.02fF
C2041 AMUX4_3V_0|SEL[0] BU_3VX2_45|Q 24.32fF
C2042 raven_padframe_0|VDDPADF_1|VDDO raven_padframe_0|VDDPADF_1|GNDO 2.28fF
C2043 BU_3VX2_37|A IN_3VX2_1|A 0.01fF
C2044 raven_padframe_0|aregc01_3v3_1|m4_0_30133# raven_padframe_0|aregc01_3v3_1|GNDR 0.07fF
C2045 raven_soc_0|gpio_in<3> BU_3VX2_63|Q 0.12fF
C2046 BU_3VX2_63|Q raven_soc_0|gpio_out<9> 0.01fF
C2047 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<12> 0.01fF
C2048 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<7> 0.01fF
C2049 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<6> 1.48fF
C2050 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<8> 0.03fF
C2051 LS_3VX2_10|A BU_3VX2_56|Q 8.77fF
C2052 LS_3VX2_24|A BU_3VX2_54|Q 0.12fF
C2053 LS_3VX2_7|A vdd 4.88fF
C2054 raven_soc_0|gpio_pulldown<4> BU_3VX2_40|Q 0.02fF
C2055 BU_3VX2_0|Q raven_soc_0|gpio_pullup<5> 0.05fF
C2056 LS_3VX2_3|A raven_soc_0|gpio_in<11> 0.53fF
C2057 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<13> 0.02fF
C2058 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<14> 0.02fF
C2059 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<9> 0.01fF
C2060 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<10> 6.51fF
C2061 raven_soc_0|gpio_pulldown<9> raven_soc_0|ext_clk 0.01fF
C2062 raven_soc_0|gpio_out<14> BU_3VX2_26|Q 0.01fF
C2063 BU_3VX2_4|Q BU_3VX2_25|Q 0.17fF
C2064 BU_3VX2_3|Q BU_3VX2_27|Q 17.23fF
C2065 BU_3VX2_32|Q apllc03_1v8_0|CLK 0.93fF
C2066 raven_soc_0|gpio_out<0> raven_soc_0|irq_pin 0.01fF
C2067 BU_3VX2_21|A BU_3VX2_19|Q 0.03fF
C2068 BU_3VX2_21|A BU_3VX2_18|Q 0.02fF
C2069 BU_3VX2_20|A raven_soc_0|flash_io1_di 0.01fF
C2070 BU_3VX2_7|A raven_soc_0|flash_clk 0.01fF
C2071 BU_3VX2_18|A raven_soc_0|flash_io0_oeb 0.01fF
C2072 BU_3VX2_40|A raven_soc_0|flash_io1_do 0.01fF
C2073 raven_soc_0|gpio_in<2> raven_soc_0|flash_io1_do 3.03fF
C2074 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<5> 0.13fF
C2075 raven_spi_0|sdo_enb raven_soc_0|flash_io2_do 0.82fF
C2076 BU_3VX2_31|A raven_soc_0|flash_io2_oeb 24.36fF
C2077 VDD raven_padframe_0|BBCUD4F_9|GNDR 0.16fF
C2078 LS_3VX2_3|A raven_soc_0|gpio_outenb<9> 0.63fF
C2079 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<6> 2.60fF
C2080 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pulldown<3> 0.01fF
C2081 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<23> 1.24fF
C2082 BU_3VX2_47|A BU_3VX2_45|A 1.28fF
C2083 BU_3VX2_47|A BU_3VX2_47|Q 0.10fF
C2084 BU_3VX2_7|A BU_3VX2_9|A 9.03fF
C2085 BU_3VX2_6|A BU_3VX2_31|A 0.01fF
C2086 BU_3VX2_23|A raven_soc_0|flash_io1_oeb 3.09fF
C2087 LS_3VX2_9|A BU_3VX2_59|Q 8.15fF
C2088 raven_soc_0|gpio_outenb<3> BU_3VX2_71|Q 0.01fF
C2089 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<10> 0.33fF
C2090 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<13> 0.30fF
C2091 raven_soc_0|gpio_in<0> BU_3VX2_28|Q 0.01fF
C2092 raven_soc_0|gpio_out<13> BU_3VX2_29|Q 0.01fF
C2093 raven_soc_0|gpio_out<11> apllc03_1v8_0|CLK 0.01fF
C2094 raven_soc_0|flash_csb BU_3VX2_28|Q 21.06fF
C2095 LS_3VX2_18|Q BU_3VX2_32|A 5.55fF
C2096 BU_3VX2_56|A BU_3VX2_56|Q 0.10fF
C2097 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<0> 12.57fF
C2098 LS_3VX2_12|A LS_3VX2_12|Q 0.05fF
C2099 VDD3V3 raven_padframe_0|VDDORPADF_3|GNDO 2.41fF
C2100 LS_3VX2_3|Q IN_3VX2_1|A 0.01fF
C2101 BU_3VX2_10|A raven_soc_0|flash_csb 0.01fF
C2102 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<14> 0.01fF
C2103 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<12> 0.01fF
C2104 BU_3VX2_33|A BU_3VX2_36|A 3.69fF
C2105 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<11> 1.78fF
C2106 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<5> 0.35fF
C2107 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<10> 19.27fF
C2108 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<12> 0.63fF
C2109 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<15> 0.02fF
C2110 BU_3VX2_0|Q raven_soc_0|gpio_outenb<12> 0.01fF
C2111 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<10> 25.18fF
C2112 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<31> 0.05fF
C2113 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<22> 0.01fF
C2114 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<30> 0.41fF
C2115 AMUX4_3V_3|SEL[1] BU_3VX2_13|Q 4.22fF
C2116 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<24> 0.03fF
C2117 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<21> 0.11fF
C2118 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<23> 0.01fF
C2119 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<10> 5.60fF
C2120 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<25> 0.42fF
C2121 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<12> 2.87fF
C2122 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<8> 28.82fF
C2123 BU_3VX2_14|Q BU_3VX2_5|Q 4.62fF
C2124 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<0> 0.04fF
C2125 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<2> 0.01fF
C2126 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<1> 0.01fF
C2127 raven_soc_0|ext_clk raven_soc_0|flash_io0_di 194.83fF
C2128 BU_3VX2_35|Q BU_3VX2_37|Q 18.69fF
C2129 BU_3VX2_40|Q raven_soc_0|flash_io2_di 13.84fF
C2130 raven_soc_0|irq_pin LS_3VX2_27|A 0.01fF
C2131 raven_soc_0|gpio_in<15> raven_padframe_0|BBCUD4F_15|PO 0.04fF
C2132 BU_3VX2_25|A BU_3VX2_16|A 2.34fF
C2133 VDD3V3 raven_padframe_0|VDDORPADF_1|GNDO 2.41fF
C2134 raven_padframe_0|ICF_1|VDDO raven_padframe_0|ICF_1|GNDO 2.28fF
C2135 BU_3VX2_25|A BU_3VX2_29|A 8.83fF
C2136 BU_3VX2_0|A raven_soc_0|flash_csb 0.01fF
C2137 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<9> 1.30fF
C2138 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<2> 3.35fF
C2139 AMUX4_3V_1|AIN1 BU_3VX2_56|A 0.02fF
C2140 BU_3VX2_68|A BU_3VX2_67|Q 0.16fF
C2141 LS_3VX2_14|A BU_3VX2_48|Q 4.71fF
C2142 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<23> 5.22fF
C2143 raven_soc_0|gpio_in<5> raven_soc_0|gpio_out<15> 0.14fF
C2144 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<28> 2.61fF
C2145 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<19> 0.01fF
C2146 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<19> 0.56fF
C2147 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<29> 0.02fF
C2148 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<25> 0.03fF
C2149 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<22> 0.04fF
C2150 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<21> 1.24fF
C2151 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<26> 0.01fF
C2152 raven_soc_0|ram_rdata<31> vdd 0.26fF
C2153 BU_3VX2_37|A BU_3VX2_25|A 0.01fF
C2154 BU_3VX2_38|A BU_3VX2_37|Q 0.03fF
C2155 BU_3VX2_6|A BU_3VX2_3|Q 0.02fF
C2156 LS_3VX2_14|A raven_soc_0|ser_tx 0.01fF
C2157 AMUX4_3V_0|AIN1 BU_3VX2_43|A 0.02fF
C2158 IN_3VX2_1|Q comp_inp 2.52fF
C2159 IN_3VX2_1|Q BU_3VX2_44|Q 1.24fF
C2160 BU_3VX2_31|A BU_3VX2_25|Q 32.45fF
C2161 raven_soc_0|gpio_pulldown<11> BU_3VX2_40|Q 0.11fF
C2162 BU_3VX2_63|Q raven_soc_0|ext_clk 42.56fF
C2163 BU_3VX2_0|Q BU_3VX2_1|Q 0.01fF
C2164 raven_soc_0|gpio_pulldown<1> BU_3VX2_26|Q 0.01fF
C2165 raven_soc_0|gpio_pulldown<2> BU_3VX2_27|Q 0.01fF
C2166 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_out<14> 33.54fF
C2167 raven_soc_0|gpio_pullup<14> BU_3VX2_71|Q 0.27fF
C2168 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<31> 16.28fF
C2169 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<10> 65.26fF
C2170 raven_padframe_0|GNDORPADF_6|VDDR raven_padframe_0|GNDORPADF_6|VDDO 0.06fF
C2171 BU_3VX2_10|A BU_3VX2_20|A 1.26fF
C2172 BU_3VX2_7|A BU_3VX2_28|A 0.01fF
C2173 LS_3VX2_14|A LS_3VX2_24|A 36.48fF
C2174 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<13> 0.01fF
C2175 BU_3VX2_3|A raven_soc_0|flash_io2_di 0.01fF
C2176 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<10> 0.01fF
C2177 BU_3VX2_22|A raven_soc_0|flash_io2_oeb 0.01fF
C2178 adc_high raven_soc_0|ser_rx 0.13fF
C2179 AMUX4_3V_4|AOUT AMUX4_3V_3|SEL[1] 0.60fF
C2180 BU_3VX2_15|A raven_soc_0|flash_io2_di 0.01fF
C2181 BU_3VX2_71|A raven_soc_0|flash_io0_oeb 0.01fF
C2182 IN_3VX2_1|A raven_soc_0|flash_io1_oeb 24.11fF
C2183 LS_3VX2_24|Q LS_3VX2_19|A 17.49fF
C2184 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<3> 0.10fF
C2185 LS_3VX2_6|A LS_3VX2_27|A 5.47fF
C2186 BU_3VX2_24|A BU_3VX2_4|A 0.01fF
C2187 acmpc01_3v3_0|IBN AMUX4_3V_3|AOUT 0.27fF
C2188 BU_3VX2_22|A BU_3VX2_6|A 0.45fF
C2189 VDD raven_padframe_0|BBC4F_1|VDDR 0.71fF
C2190 VDD raven_padframe_0|ICF_1|VDDR 0.71fF
C2191 BU_3VX2_20|A BU_3VX2_0|A 0.01fF
C2192 raven_soc_0|gpio_pullup<2> LS_3VX2_3|A 0.01fF
C2193 BU_3VX2_31|A BU_3VX2_27|A 13.55fF
C2194 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<1> 21.32fF
C2195 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<4> 5.80fF
C2196 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<15> 0.21fF
C2197 raven_soc_0|gpio_out<11> raven_soc_0|gpio_outenb<8> 0.02fF
C2198 raven_soc_0|gpio_in<0> raven_padframe_0|BBCUD4F_1|PO 0.04fF
C2199 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<27> 2.70fF
C2200 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<21> 0.01fF
C2201 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<7> 4.19fF
C2202 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<6> 5.39fF
C2203 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<27> 4.06fF
C2204 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<25> 9.83fF
C2205 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<22> 2.85fF
C2206 LS_3VX2_2|A BU_3VX2_33|Q 27.39fF
C2207 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<21> 20.31fF
C2208 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<15> 16.97fF
C2209 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<17> 0.11fF
C2210 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<1> 0.04fF
C2211 raven_soc_0|gpio_in<10> vdd 2.21fF
C2212 raven_soc_0|gpio_in<12> apllc03_1v8_0|CLK 0.06fF
C2213 raven_soc_0|gpio_in<14> BU_3VX2_29|Q 0.01fF
C2214 raven_soc_0|ser_tx BU_3VX2_56|Q 6.06fF
C2215 VDD3V3 BU_3VX2_62|Q 0.05fF
C2216 raven_soc_0|gpio_in<13> BU_3VX2_28|Q 0.01fF
C2217 BU_3VX2_42|Q BU_3VX2_72|Q 5.58fF
C2218 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<14> 0.01fF
C2219 BU_3VX2_25|A LS_3VX2_3|Q 0.01fF
C2220 raven_padframe_0|ICF_1|VDDR LOGIC0_3V_4|Q 0.01fF
C2221 raven_padframe_0|BBC4F_1|VDDR LOGIC0_3V_4|Q 0.01fF
C2222 AMUX4_3V_0|AIN1 adc_low 0.27fF
C2223 LOGIC1_3V_1|Q LOGIC0_3V_2|Q 2.89fF
C2224 LS_3VX2_9|A AMUX2_3V_0|SEL 8.83fF
C2225 raven_padframe_0|aregc01_3v3_1|m4_92500_30133# raven_padframe_0|aregc01_3v3_1|m4_92500_29333# 0.09fF
C2226 raven_padframe_0|aregc01_3v3_1|m4_0_29057# raven_padframe_0|aregc01_3v3_1|m4_0_22024# 0.02fF
C2227 raven_padframe_0|aregc01_3v3_1|m4_92500_30653# raven_padframe_0|aregc01_3v3_1|m4_92500_29057# 0.01fF
C2228 LS_3VX2_10|Q LS_3VX2_6|A 0.54fF
C2229 adc_low LS_3VX2_24|Q 3.52fF
C2230 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<7> 0.01fF
C2231 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<8> 98.89fF
C2232 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<4> 0.22fF
C2233 BU_3VX2_63|Q raven_soc_0|gpio_outenb<10> 0.01fF
C2234 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<5> 0.01fF
C2235 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<12> 0.01fF
C2236 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<7> 0.17fF
C2237 LS_3VX2_5|A VDD3V3 0.52fF
C2238 LS_3VX2_24|A BU_3VX2_56|Q 0.02fF
C2239 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<13> 28.14fF
C2240 BU_3VX2_1|Q raven_soc_0|flash_io3_di 0.01fF
C2241 BU_3VX2_3|Q BU_3VX2_25|Q 3.90fF
C2242 BU_3VX2_14|Q BU_3VX2_28|Q 0.03fF
C2243 BU_3VX2_37|Q BU_3VX2_23|Q 0.01fF
C2244 raven_soc_0|gpio_out<10> BU_3VX2_24|Q 0.01fF
C2245 LS_3VX2_22|A adc0_data<5> 4.76fF
C2246 raven_soc_0|ram_rdata<16> apllc03_1v8_0|CLK 0.01fF
C2247 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<3> 8.52fF
C2248 BU_3VX2_16|A BU_3VX2_13|Q 0.02fF
C2249 BU_3VX2_5|A raven_soc_0|ext_clk 0.04fF
C2250 BU_3VX2_18|A raven_soc_0|flash_io2_do 0.01fF
C2251 LS_3VX2_6|Q LS_3VX2_19|A 0.01fF
C2252 IN_3VX2_1|Q vdd 0.12fF
C2253 raven_padframe_0|BBC4F_1|VDDR raven_padframe_0|BBC4F_1|VDDO 0.06fF
C2254 raven_padframe_0|BT4F_2|VDDR raven_padframe_0|BT4F_2|GNDR 0.68fF
C2255 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<10> 6.68fF
C2256 analog_out AMUX4_3V_4|AIN3 6.99fF
C2257 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<3> 0.16fF
C2258 BU_3VX2_0|Q raven_soc_0|ram_wdata<29> 0.02fF
C2259 raven_soc_0|gpio_outenb<2> VDD3V3 2.48fF
C2260 raven_soc_0|gpio_out<2> raven_soc_0|ext_clk 0.01fF
C2261 BU_3VX2_51|A BU_3VX2_41|A 0.96fF
C2262 BU_3VX2_49|A BU_3VX2_48|A 11.16fF
C2263 BU_3VX2_50|A BU_3VX2_47|A 1.94fF
C2264 raven_padframe_0|APR00DF_4|GNDR raven_padframe_0|APR00DF_4|VDDO 0.09fF
C2265 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<13> 1.24fF
C2266 BU_3VX2_21|A raven_soc_0|flash_io2_oeb 0.01fF
C2267 LS_3VX2_8|Q LS_3VX2_19|A 0.01fF
C2268 LS_3VX2_9|A BU_3VX2_61|Q 6.51fF
C2269 raven_soc_0|gpio_out<0> BU_3VX2_26|Q 0.01fF
C2270 BU_3VX2_17|A raven_soc_0|flash_io3_oeb 0.01fF
C2271 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<14> 0.97fF
C2272 aopac01_3v3_0|IB vdd 0.01fF
C2273 raven_soc_0|gpio_in<0> vdd 3.43fF
C2274 raven_soc_0|flash_csb vdd 0.16fF
C2275 raven_soc_0|gpio_outenb<15> BU_3VX2_29|Q 0.01fF
C2276 raven_soc_0|gpio_out<12> BU_3VX2_26|Q 0.01fF
C2277 raven_soc_0|gpio_outenb<11> BU_3VX2_27|Q 0.01fF
C2278 BU_3VX2_35|Q BU_3VX2_40|Q 0.45fF
C2279 BU_3VX2_6|A BU_3VX2_21|A 0.58fF
C2280 VDD raven_padframe_0|GNDORPADF_5|VDDR 0.71fF
C2281 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<10> 0.01fF
C2282 LS_3VX2_13|Q LS_3VX2_14|Q 0.28fF
C2283 BU_3VX2_4|A BU_3VX2_16|A 0.85fF
C2284 BU_3VX2_7|A BU_3VX2_14|A 1.66fF
C2285 BU_3VX2_4|A BU_3VX2_29|A 0.01fF
C2286 LS_3VX2_6|Q adc_low 0.12fF
C2287 IN_3VX2_1|A raven_soc_0|gpio_pulldown<13> 0.01fF
C2288 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<7> 0.62fF
C2289 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<9> 0.08fF
C2290 LS_3VX2_3|A raven_soc_0|gpio_outenb<14> 0.01fF
C2291 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<5> 0.01fF
C2292 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<10> 12.15fF
C2293 BU_3VX2_25|A raven_soc_0|flash_io1_oeb 3.28fF
C2294 BU_3VX2_0|Q raven_soc_0|gpio_pullup<12> 0.01fF
C2295 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<7> 0.01fF
C2296 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<30> 0.20fF
C2297 raven_soc_0|ram_wenb raven_soc_0|ram_addr<2> 0.01fF
C2298 raven_soc_0|gpio_in<11> raven_soc_0|gpio_in<10> 25.28fF
C2299 AMUX4_3V_3|SEL[1] BU_3VX2_69|Q 1.52fF
C2300 raven_soc_0|gpio_in<6> raven_soc_0|gpio_out<15> 0.09fF
C2301 VDD3V3 BU_3VX2_45|Q 1.52fF
C2302 VDD raven_padframe_0|BBCUD4F_14|VDDR 0.71fF
C2303 raven_padframe_0|GNDORPADF_5|VDDR LOGIC0_3V_4|Q 0.01fF
C2304 BU_3VX2_37|A BU_3VX2_4|A 3.15fF
C2305 LS_3VX2_8|Q adc_low 0.12fF
C2306 BU_3VX2_22|A BU_3VX2_27|A 4.45fF
C2307 BU_3VX2_40|A raven_soc_0|flash_csb 0.01fF
C2308 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<2> 9.56fF
C2309 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<3> 0.01fF
C2310 IN_3VX2_1|A raven_soc_0|gpio_pullup<1> 0.01fF
C2311 raven_padframe_0|aregc01_3v3_0|m4_0_30653# raven_padframe_0|aregc01_3v3_0|VDDR 0.07fF
C2312 raven_padframe_0|aregc01_3v3_0|m4_92500_30133# raven_padframe_0|aregc01_3v3_0|m4_92500_29057# 0.01fF
C2313 LS_3VX2_24|Q AMUX2_3V_0|AOUT 0.01fF
C2314 LOGIC0_3V_3|Q BU_3VX2_33|A 1.17fF
C2315 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<6> 1.05fF
C2316 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<10> 0.36fF
C2317 BU_3VX2_68|A BU_3VX2_65|Q 0.02fF
C2318 BU_3VX2_38|A BU_3VX2_40|Q 0.03fF
C2319 BU_3VX2_71|Q raven_soc_0|gpio_in<9> 0.06fF
C2320 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<19> 0.04fF
C2321 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<6> 10.63fF
C2322 raven_soc_0|gpio_out<10> raven_soc_0|gpio_out<15> 0.64fF
C2323 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<28> 171.29fF
C2324 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<10> 9.27fF
C2325 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<20> 13.50fF
C2326 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<11> 0.01fF
C2327 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<0> 5.95fF
C2328 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<23> 0.09fF
C2329 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<12> 0.02fF
C2330 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<8> 0.01fF
C2331 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<13> 0.02fF
C2332 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<14> 0.01fF
C2333 raven_soc_0|ram_rdata<30> vdd 0.30fF
C2334 raven_soc_0|ram_rdata<22> apllc03_1v8_0|CLK 0.01fF
C2335 AMUX4_3V_0|SEL[0] LS_3VX2_21|A 0.01fF
C2336 BU_3VX2_20|A vdd 0.06fF
C2337 LS_3VX2_8|A LS_3VX2_20|A 5.78fF
C2338 BU_3VX2_12|A raven_soc_0|flash_io3_oeb 0.01fF
C2339 BU_3VX2_26|A raven_soc_0|flash_io3_do 0.01fF
C2340 VDD raven_padframe_0|APR00DF_2|GNDR 0.16fF
C2341 raven_soc_0|gpio_outenb<1> BU_3VX2_28|Q 0.01fF
C2342 raven_soc_0|gpio_pulldown<2> BU_3VX2_25|Q 0.01fF
C2343 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<31> 12.66fF
C2344 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<6> 1.41fF
C2345 raven_soc_0|ram_addr<4> raven_soc_0|ram_addr<2> 33.92fF
C2346 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<7> 6.39fF
C2347 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<10> 11.68fF
C2348 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<24> 1.98fF
C2349 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<5> 0.03fF
C2350 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_out<14> 206.61fF
C2351 BU_3VX2_37|Q BU_3VX2_4|Q 14.58fF
C2352 raven_soc_0|gpio_in<1> raven_soc_0|flash_io1_di 0.46fF
C2353 BU_3VX2_2|A BU_3VX2_12|A 1.50fF
C2354 BU_3VX2_24|A raven_soc_0|flash_io0_oeb 3.61fF
C2355 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<12> 0.01fF
C2356 BU_3VX2_71|A raven_soc_0|flash_io2_do 0.01fF
C2357 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<7> 0.01fF
C2358 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<11> 4.61fF
C2359 LS_3VX2_24|Q LS_3VX2_22|A 8.80fF
C2360 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<15> 0.01fF
C2361 BU_3VX2_11|A raven_soc_0|flash_io3_do 0.01fF
C2362 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<15> 1.06fF
C2363 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<15> 0.56fF
C2364 LOGIC0_3V_1|Q raven_spi_0|SDO 2.83fF
C2365 BU_3VX2_3|A BU_3VX2_38|A 3.00fF
C2366 BU_3VX2_4|A LS_3VX2_3|Q 0.49fF
C2367 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<13> 0.34fF
C2368 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<9> 0.01fF
C2369 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<5> 1.18fF
C2370 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<5> 0.71fF
C2371 raven_soc_0|gpio_out<12> raven_soc_0|gpio_outenb<13> 16.76fF
C2372 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<2> 4.53fF
C2373 BU_3VX2_15|Q BU_3VX2_21|Q 5.68fF
C2374 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<22> 13.33fF
C2375 BU_3VX2_38|Q BU_3VX2_13|Q 2.69fF
C2376 raven_soc_0|ram_rdata<3> raven_soc_0|ram_addr<1> 0.30fF
C2377 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<26> 2.39fF
C2378 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<1> 0.01fF
C2379 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<25> 3.67fF
C2380 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<21> 12.45fF
C2381 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<25> 11.46fF
C2382 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<8> 0.01fF
C2383 BU_3VX2_22|Q BU_3VX2_10|Q 2.88fF
C2384 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<17> 23.17fF
C2385 BU_3VX2_15|Q BU_3VX2_8|Q 5.00fF
C2386 BU_3VX2_13|Q BU_3VX2_67|Q 7.10fF
C2387 BU_3VX2_21|Q BU_3VX2_9|Q 11.56fF
C2388 BU_3VX2_2|Q BU_3VX2_22|Q 0.05fF
C2389 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<19> 16.16fF
C2390 BU_3VX2_1|Q AMUX4_3V_3|SEL[0] 0.86fF
C2391 BU_3VX2_12|Q BU_3VX2_20|Q 4.07fF
C2392 BU_3VX2_9|Q BU_3VX2_8|Q 68.01fF
C2393 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<26> 6.24fF
C2394 BU_3VX2_6|Q BU_3VX2_17|Q 2.92fF
C2395 BU_3VX2_7|Q BU_3VX2_17|Q 3.31fF
C2396 raven_soc_0|gpio_in<13> vdd 1.40fF
C2397 raven_soc_0|ext_clk BU_3VX2_24|Q 0.01fF
C2398 BU_3VX2_40|Q BU_3VX2_23|Q 0.01fF
C2399 BU_3VX2_59|A vdd 0.17fF
C2400 raven_padframe_0|FILLER50F_2|VDDO raven_padframe_0|FILLER50F_2|GNDO 2.28fF
C2401 raven_padframe_0|BBC4F_1|GNDR raven_padframe_0|BBC4F_1|GNDO 0.81fF
C2402 raven_padframe_0|FILLER20F_7|VDDO raven_padframe_0|FILLER20F_7|GNDO 2.28fF
C2403 BU_3VX2_21|A BU_3VX2_27|A 3.58fF
C2404 raven_padframe_0|aregc01_3v3_1|m4_0_29333# raven_padframe_0|aregc01_3v3_1|m4_0_29057# 0.11fF
C2405 raven_padframe_0|aregc01_3v3_1|m4_0_30133# raven_padframe_0|aregc01_3v3_1|m4_0_28769# 0.01fF
C2406 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<9> 7.97fF
C2407 raven_padframe_0|axtoc02_3v3_0|m4_0_30653# raven_padframe_0|axtoc02_3v3_0|m4_0_29333# 0.03fF
C2408 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<7> 0.01fF
C2409 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<0> 0.01fF
C2410 BU_3VX2_63|Q raven_soc_0|gpio_pullup<10> 0.01fF
C2411 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<6> 0.01fF
C2412 raven_soc_0|gpio_out<4> BU_3VX2_40|Q 0.11fF
C2413 AMUX4_3V_3|SEL[1] BU_3VX2_29|Q 0.05fF
C2414 BU_3VX2_14|Q vdd 2.35fF
C2415 raven_soc_0|gpio_pulldown<7> apllc03_1v8_0|CLK 0.43fF
C2416 BU_3VX2_35|A LOGIC0_3V_2|Q 0.06fF
C2417 raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<11> 10.61fF
C2418 markings_0|product_name_0|_alphabet_E_0|m2_0_0# markings_0|product_name_0|_alphabet_A_0|m2_0_0# 0.12fF
C2419 markings_0|manufacturer_0|_alphabet_E_1|m2_0_0# markings_0|product_name_0|_alphabet_R_0|m2_0_0# 0.15fF
C2420 BU_3VX2_7|A raven_soc_0|flash_io1_do 0.01fF
C2421 acsoc01_3v3_0|CS3_200N VDD3V3 0.02fF
C2422 acsoc02_3v3_0|CS_4U VDD3V3 0.02fF
C2423 LS_3VX2_6|Q LS_3VX2_22|A 0.01fF
C2424 BU_3VX2_31|A raven_soc_0|gpio_in<7> 0.01fF
C2425 BU_3VX2_13|A raven_soc_0|ext_clk 0.01fF
C2426 VDD raven_padframe_0|FILLER20F_6|GNDO 0.07fF
C2427 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<3> 0.57fF
C2428 AMUX4_3V_4|AIN1 AMUX4_3V_4|AIN3 24.65fF
C2429 BU_3VX2_0|Q raven_soc_0|ram_rdata<29> 3.18fF
C2430 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<13> 0.01fF
C2431 BU_3VX2_33|A VDD3V3 1.32fF
C2432 raven_soc_0|flash_io2_di raven_soc_0|ram_rdata<11> 0.05fF
C2433 raven_soc_0|ram_rdata<10> raven_soc_0|ram_addr<0> 0.09fF
C2434 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<15> 0.83fF
C2435 BU_3VX2_48|A BU_3VX2_46|Q 0.02fF
C2436 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<15> 0.89fF
C2437 raven_padframe_0|FILLER10F_0|VDDO raven_padframe_0|FILLER10F_0|GNDO 2.28fF
C2438 raven_soc_0|gpio_in<1> BU_3VX2_28|Q 0.01fF
C2439 LS_3VX2_9|A LS_3VX2_15|A 0.02fF
C2440 LS_3VX2_8|Q LS_3VX2_22|A 0.01fF
C2441 LS_3VX2_12|A BU_3VX2_55|Q 6.25fF
C2442 BU_3VX2_4|A raven_soc_0|flash_io1_oeb 0.01fF
C2443 BU_3VX2_16|A raven_soc_0|flash_io0_oeb 0.01fF
C2444 VDD raven_padframe_0|BBC4F_0|GNDR 0.16fF
C2445 raven_soc_0|gpio_pullup<0> BU_3VX2_71|Q 0.01fF
C2446 BU_3VX2_29|A raven_soc_0|flash_io0_oeb 9.95fF
C2447 IN_3VX2_1|A BU_3VX2_72|Q 7.17fF
C2448 raven_soc_0|gpio_pullup<11> BU_3VX2_27|Q 0.01fF
C2449 raven_soc_0|gpio_outenb<10> BU_3VX2_24|Q 0.01fF
C2450 LS_3VX2_13|A BU_3VX2_54|Q 0.01fF
C2451 raven_soc_0|gpio_outenb<12> BU_3VX2_26|Q 0.01fF
C2452 raven_soc_0|gpio_outenb<11> BU_3VX2_25|Q 0.01fF
C2453 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<12> 0.01fF
C2454 LS_3VX2_13|Q LS_3VX2_7|Q 3.10fF
C2455 BU_3VX2_8|A BU_3VX2_26|A 0.01fF
C2456 BU_3VX2_1|A BU_3VX2_36|A 0.67fF
C2457 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<7> 1.93fF
C2458 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<3> 0.01fF
C2459 BU_3VX2_37|A raven_soc_0|flash_io0_oeb 0.01fF
C2460 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<7> 0.02fF
C2461 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pulldown<4> 0.46fF
C2462 LS_3VX2_3|A raven_soc_0|gpio_pullup<15> 0.01fF
C2463 BU_3VX2_35|A raven_soc_0|flash_io0_do 0.07fF
C2464 BU_3VX2_0|Q raven_soc_0|gpio_outenb<0> 0.01fF
C2465 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<5> 0.01fF
C2466 AMUX4_3V_4|AOUT raven_soc_0|flash_io1_oeb 1.88fF
C2467 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<8> 0.10fF
C2468 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<11> 24.00fF
C2469 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<15> 2.09fF
C2470 raven_soc_0|ext_clk raven_soc_0|gpio_out<15> 0.01fF
C2471 raven_soc_0|flash_io3_do VDD3V3 10.60fF
C2472 VDD3V3 AMUX4_3V_4|AIN3 17.34fF
C2473 BU_3VX2_60|A LS_3VX2_17|Q 0.29fF
C2474 BU_3VX2_59|A BU_3VX2_62|A 0.28fF
C2475 BU_3VX2_61|A LS_3VX2_16|Q 1.21fF
C2476 AMUX4_3V_1|AOUT comp_inp 1.20fF
C2477 raven_soc_0|irq_pin BU_3VX2_53|Q 0.01fF
C2478 LS_3VX2_20|A BU_3VX2_44|Q 10.18fF
C2479 raven_padframe_0|FILLER20FC_0|VDDO raven_padframe_0|FILLER20FC_0|GNDO 2.28fF
C2480 BU_3VX2_8|A BU_3VX2_11|A 4.41fF
C2481 raven_padframe_0|APR00DF_5|GNDR raven_padframe_0|APR00DF_5|GNDO 0.81fF
C2482 raven_padframe_0|FILLER20F_4|VDDR raven_padframe_0|FILLER20F_4|GNDO 0.13fF
C2483 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_outenb<0> 49.09fF
C2484 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<5> 0.01fF
C2485 BU_3VX2_31|A raven_soc_0|gpio_out<7> 0.01fF
C2486 raven_padframe_0|aregc01_3v3_0|m4_0_29333# raven_padframe_0|aregc01_3v3_0|m4_0_28769# 0.03fF
C2487 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<3> 2.18fF
C2488 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<10> 0.01fF
C2489 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<8> 0.02fF
C2490 markings_0|efabless_logo_0|m1_2700_n10050# markings_0|efabless_logo_0|m1_3600_n10650# 0.33fF
C2491 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<13> 0.02fF
C2492 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<6> 0.12fF
C2493 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<20> 0.01fF
C2494 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<7> 11.29fF
C2495 raven_soc_0|gpio_in<5> raven_soc_0|ext_clk 0.01fF
C2496 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<0> 0.01fF
C2497 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_pullup<5> 0.02fF
C2498 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<9> 0.01fF
C2499 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<12> 6.63fF
C2500 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<25> 36.10fF
C2501 raven_soc_0|gpio_out<14> VDD3V3 0.07fF
C2502 BU_3VX2_73|Q BU_3VX2_59|Q 0.01fF
C2503 raven_soc_0|ram_rdata<7> vdd 0.36fF
C2504 AMUX4_3V_0|SEL[0] LS_3VX2_27|A 0.01fF
C2505 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_in<0> 4.36fF
C2506 raven_padframe_0|VDDPADF_0|VDDR raven_padframe_0|VDDPADF_0|GNDR 0.68fF
C2507 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<6> 5.75fF
C2508 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<15> 37.23fF
C2509 LS_3VX2_11|A VDD3V3 0.51fF
C2510 VDD raven_padframe_0|CORNERESDF_3|VDDR 0.71fF
C2511 VDD raven_padframe_0|BBCUD4F_7|GNDO 0.07fF
C2512 BU_3VX2_0|Q BU_3VX2_12|Q 0.01fF
C2513 raven_soc_0|gpio_outenb<1> vdd 0.19fF
C2514 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_outenb<8> 14.79fF
C2515 raven_soc_0|ram_rdata<14> raven_soc_0|ram_addr<3> 0.44fF
C2516 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<7> 0.05fF
C2517 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<9> 0.95fF
C2518 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<30> 15.29fF
C2519 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<8> 6.92fF
C2520 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<6> 52.03fF
C2521 raven_soc_0|ram_rdata<5> raven_soc_0|ram_addr<2> 0.31fF
C2522 raven_soc_0|ram_rdata<18> raven_soc_0|ram_addr<4> 0.01fF
C2523 BU_3VX2_37|Q BU_3VX2_3|Q 24.95fF
C2524 BU_3VX2_14|Q BU_3VX2_70|Q 3.04fF
C2525 raven_soc_0|ram_rdata<23> apllc03_1v8_0|CLK 0.01fF
C2526 raven_padframe_0|APR00DF_1|GNDR raven_padframe_0|APR00DF_1|VDDO 0.09fF
C2527 raven_padframe_0|axtoc02_3v3_0|VDDR raven_padframe_0|axtoc02_3v3_0|GNDR 0.93fF
C2528 BU_3VX2_24|A raven_soc_0|flash_io2_do 0.01fF
C2529 LS_3VX2_9|A AMUX4_3V_1|SEL[1] 63.87fF
C2530 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<8> 1.17fF
C2531 LS_3VX2_14|Q LS_3VX2_19|A 0.36fF
C2532 LS_3VX2_3|Q raven_soc_0|flash_io0_oeb 0.01fF
C2533 IN_3VX2_1|A AMUX4_3V_1|SEL[0] 0.01fF
C2534 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<6> 0.87fF
C2535 LS_3VX2_6|A BU_3VX2_53|Q 10.97fF
C2536 BU_3VX2_29|A BU_3VX2_29|Q 0.08fF
C2537 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<10> 0.19fF
C2538 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<14> 0.64fF
C2539 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<12> 38.43fF
C2540 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<6> 1.73fF
C2541 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<7> 1.54fF
C2542 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<8> 1.05fF
C2543 BU_3VX2_0|Q raven_soc_0|flash_io0_do 0.01fF
C2544 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<15> 0.02fF
C2545 raven_padframe_0|APR00DF_1|VDDR raven_padframe_0|APR00DF_1|VDDO 0.06fF
C2546 LS_3VX2_9|A LS_3VX2_7|A 17.99fF
C2547 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<3> 2.01fF
C2548 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<13> 0.01fF
C2549 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_in<2> 10.36fF
C2550 BU_3VX2_3|A BU_3VX2_4|Q 0.03fF
C2551 LOGIC0_3V_4|Q raven_soc_0|flash_io0_oeb 0.01fF
C2552 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<10> 0.01fF
C2553 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<8> 15.55fF
C2554 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<10> 23.35fF
C2555 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<13> 26.81fF
C2556 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<5> 0.01fF
C2557 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pullup<6> 0.02fF
C2558 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pullup<13> 10.88fF
C2559 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<14> 0.02fF
C2560 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<13> 0.78fF
C2561 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<1> 0.01fF
C2562 raven_soc_0|gpio_pulldown<8> BU_3VX2_27|Q 0.01fF
C2563 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<26> 2.58fF
C2564 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<27> 0.84fF
C2565 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<3> 3.69fF
C2566 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<2> 0.01fF
C2567 BU_3VX2_66|Q BU_3VX2_5|Q 1.24fF
C2568 BU_3VX2_16|Q BU_3VX2_12|Q 12.83fF
C2569 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<13> 9.28fF
C2570 BU_3VX2_19|Q BU_3VX2_9|Q 3.26fF
C2571 BU_3VX2_21|Q BU_3VX2_64|Q 1.00fF
C2572 BU_3VX2_38|Q BU_3VX2_69|Q 0.59fF
C2573 BU_3VX2_13|Q BU_3VX2_65|Q 11.99fF
C2574 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<13> 11.59fF
C2575 BU_3VX2_12|Q BU_3VX2_30|Q 2.92fF
C2576 BU_3VX2_19|Q BU_3VX2_15|Q 9.23fF
C2577 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<8> 0.18fF
C2578 BU_3VX2_35|Q BU_3VX2_17|Q 0.01fF
C2579 BU_3VX2_15|Q BU_3VX2_18|Q 13.01fF
C2580 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<17> 11.30fF
C2581 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<19> 4.05fF
C2582 BU_3VX2_69|Q BU_3VX2_67|Q 11.12fF
C2583 BU_3VX2_64|Q BU_3VX2_8|Q 0.01fF
C2584 BU_3VX2_18|Q BU_3VX2_9|Q 4.21fF
C2585 BU_3VX2_31|Q BU_3VX2_10|Q 6.62fF
C2586 LS_3VX2_20|A vdd 3.03fF
C2587 raven_padframe_0|FILLER20F_6|VDDO raven_padframe_0|FILLER20F_6|GNDO 2.28fF
C2588 LS_3VX2_14|A LS_3VX2_13|A 150.65fF
C2589 LS_3VX2_14|Q adc_low 0.33fF
C2590 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<2> 0.16fF
C2591 raven_soc_0|gpio_out<3> LS_3VX2_3|A 0.01fF
C2592 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<4> 0.71fF
C2593 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<10> 0.81fF
C2594 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<9> 9.44fF
C2595 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<4> 0.01fF
C2596 raven_soc_0|gpio_pulldown<14> BU_3VX2_0|Q 0.01fF
C2597 raven_soc_0|gpio_pulldown<3> vdd 0.15fF
C2598 raven_soc_0|ram_rdata<1> vdd 0.70fF
C2599 VDD3V3 LS_3VX2_21|A 0.50fF
C2600 raven_soc_0|ram_wdata<21> apllc03_1v8_0|CLK 0.01fF
C2601 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<5> 0.21fF
C2602 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<14> 0.42fF
C2603 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<9> 0.01fF
C2604 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<14> 0.01fF
C2605 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<6> 6.11fF
C2606 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<11> 0.01fF
C2607 markings_0|product_name_0|_alphabet_N_0|m2_0_0# markings_0|product_name_0|_alphabet_V_0|m2_0_560# 0.13fF
C2608 markings_0|efabless_logo_0|m1_3300_n1350# markings_0|efabless_logo_0|m1_7500_n3450# 0.01fF
C2609 BU_3VX2_2|A BU_3VX2_2|Q 0.08fF
C2610 BU_3VX2_8|A VDD3V3 0.19fF
C2611 raven_soc_0|gpio_pulldown<1> VDD3V3 1.81fF
C2612 BU_3VX2_0|Q raven_soc_0|ram_rdata<25> 0.02fF
C2613 raven_soc_0|flash_io3_oeb raven_soc_0|flash_clk 52.42fF
C2614 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<29> 2.97fF
C2615 raven_soc_0|flash_io0_di raven_soc_0|flash_io2_di 181.20fF
C2616 raven_soc_0|flash_io3_di raven_soc_0|flash_io0_do 60.12fF
C2617 raven_soc_0|flash_io0_oeb raven_soc_0|flash_io1_oeb 382.25fF
C2618 raven_soc_0|ram_addr<3> raven_soc_0|ram_addr<0> 20.56fF
C2619 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<1> 3.85fF
C2620 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<15> 5.01fF
C2621 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<13> 0.62fF
C2622 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<17> 0.01fF
C2623 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<16> 1.75fF
C2624 BU_3VX2_45|A BU_3VX2_44|Q 0.14fF
C2625 BU_3VX2_45|Q adc0_data<5> 75.66fF
C2626 BU_3VX2_44|Q BU_3VX2_47|Q 33.03fF
C2627 raven_padframe_0|ICFC_0|GNDR raven_padframe_0|ICFC_0|GNDO 0.81fF
C2628 raven_padframe_0|GNDORPADF_0|VDDO raven_padframe_0|GNDORPADF_0|GNDOR 2.38fF
C2629 raven_padframe_0|VDDORPADF_1|GNDR raven_padframe_0|VDDORPADF_1|GNDO 0.81fF
C2630 raven_padframe_0|FILLER20F_3|GNDR raven_padframe_0|FILLER20F_3|VDDO 0.09fF
C2631 raven_soc_0|gpio_in<1> vdd 1.34fF
C2632 BU_3VX2_9|A raven_soc_0|flash_io3_oeb 0.01fF
C2633 BU_3VX2_2|A raven_soc_0|flash_clk 0.01fF
C2634 VDD BU_3VX2_29|Q 0.05fF
C2635 BU_3VX2_16|A raven_soc_0|flash_io2_do 0.06fF
C2636 LS_3VX2_12|A BU_3VX2_57|Q 0.01fF
C2637 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<14> 0.81fF
C2638 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<9> 0.51fF
C2639 BU_3VX2_29|A raven_soc_0|flash_io2_do 4.15fF
C2640 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<3> 1.96fF
C2641 BU_3VX2_36|A BU_3VX2_1|Q 0.16fF
C2642 AMUX2_3V_0|SEL BU_3VX2_73|Q 48.85fF
C2643 IN_3VX2_1|A LS_3VX2_17|A 0.01fF
C2644 LS_3VX2_13|A BU_3VX2_56|Q 3.48fF
C2645 raven_soc_0|gpio_outenb<5> vdd 0.19fF
C2646 raven_soc_0|gpio_pullup<9> BU_3VX2_23|Q 0.01fF
C2647 raven_soc_0|gpio_pullup<11> BU_3VX2_25|Q 0.01fF
C2648 raven_soc_0|gpio_pullup<4> apllc03_1v8_0|CLK 0.01fF
C2649 raven_soc_0|gpio_pullup<12> BU_3VX2_26|Q 0.01fF
C2650 raven_soc_0|gpio_pullup<7> BU_3VX2_28|Q 0.01fF
C2651 raven_soc_0|gpio_pullup<10> BU_3VX2_24|Q 0.01fF
C2652 BU_3VX2_2|A BU_3VX2_9|A 1.17fF
C2653 LS_3VX2_13|Q LS_3VX2_4|Q 0.40fF
C2654 LS_3VX2_14|A raven_soc_0|ser_rx 0.01fF
C2655 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<5> 0.98fF
C2656 BU_3VX2_37|A raven_soc_0|flash_io2_do 0.01fF
C2657 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<9> 0.01fF
C2658 BU_3VX2_35|A raven_soc_0|flash_io1_di 0.12fF
C2659 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<7> 0.01fF
C2660 raven_soc_0|gpio_pulldown<10> BU_3VX2_0|Q 0.01fF
C2661 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<6> 1.24fF
C2662 BU_3VX2_63|Q raven_soc_0|flash_io2_di 11.43fF
C2663 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<12> 24.56fF
C2664 raven_soc_0|ext_clk raven_soc_0|gpio_in<6> 0.01fF
C2665 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<8> 0.44fF
C2666 BU_3VX2_56|A BU_3VX2_58|A 2.92fF
C2667 BU_3VX2_53|A BU_3VX2_61|A 0.28fF
C2668 BU_3VX2_52|A LS_3VX2_15|Q 0.13fF
C2669 BU_3VX2_54|A BU_3VX2_60|A 0.48fF
C2670 BU_3VX2_55|A BU_3VX2_59|A 0.92fF
C2671 VDD3V3 LS_3VX2_17|Q 1.28fF
C2672 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<2> 16.54fF
C2673 raven_padframe_0|ICFC_0|VDDR raven_padframe_0|ICFC_0|VDD3 0.71fF
C2674 raven_soc_0|gpio_in<13> raven_padframe_0|BBCUD4F_13|PO 0.04fF
C2675 BU_3VX2_3|A BU_3VX2_31|A 0.01fF
C2676 BU_3VX2_15|A BU_3VX2_31|A 0.01fF
C2677 BU_3VX2_7|A raven_soc_0|flash_csb 0.01fF
C2678 BU_3VX2_67|A BU_3VX2_70|A 4.89fF
C2679 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<10> 0.32fF
C2680 BU_3VX2_31|A raven_soc_0|gpio_outenb<7> 0.01fF
C2681 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<5> 0.01fF
C2682 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<4> 0.25fF
C2683 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<5> 0.01fF
C2684 markings_0|efabless_logo_0|m1_600_n4050# markings_0|efabless_logo_0|m1_0_n4950# 0.22fF
C2685 LOGIC0_3V_0|Q LOGIC1_3V_1|Q 0.21fF
C2686 raven_soc_0|gpio_out<8> BU_3VX2_40|Q 0.16fF
C2687 raven_soc_0|flash_io0_do raven_soc_0|irq_pin 0.07fF
C2688 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_pullup<5> 0.03fF
C2689 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<12> 0.02fF
C2690 raven_soc_0|gpio_out<10> raven_soc_0|ext_clk 0.01fF
C2691 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<7> 5.09fF
C2692 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<15> 0.02fF
C2693 raven_soc_0|ser_tx AMUX4_3V_4|AIN2 9.89fF
C2694 BU_3VX2_66|Q BU_3VX2_28|Q 0.05fF
C2695 BU_3VX2_38|Q BU_3VX2_29|Q 0.01fF
C2696 BU_3VX2_15|Q BU_3VX2_27|Q 2.93fF
C2697 BU_3VX2_73|Q BU_3VX2_61|Q 0.01fF
C2698 BU_3VX2_2|Q apllc03_1v8_0|CLK 0.01fF
C2699 BU_3VX2_17|Q BU_3VX2_23|Q 8.75fF
C2700 BU_3VX2_67|Q BU_3VX2_29|Q 0.91fF
C2701 BU_3VX2_9|Q BU_3VX2_27|Q 0.02fF
C2702 BU_3VX2_20|Q BU_3VX2_28|Q 4.25fF
C2703 BU_3VX2_10|Q apllc03_1v8_0|CLK 0.01fF
C2704 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<11> 0.01fF
C2705 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<11> 0.01fF
C2706 raven_padframe_0|FILLER20FC_0|VDDR raven_padframe_0|FILLER20FC_0|GNDR 0.68fF
C2707 LS_3VX2_24|A AMUX4_3V_4|AIN2 2.00fF
C2708 raven_soc_0|ser_rx BU_3VX2_56|Q 1.83fF
C2709 BU_3VX2_0|Q BU_3VX2_5|Q 0.01fF
C2710 raven_soc_0|ram_rdata<15> raven_soc_0|ram_rdata<16> 91.02fF
C2711 AMUX4_3V_3|SEL[1] BU_3VX2_32|Q 6.75fF
C2712 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<24> 0.08fF
C2713 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<18> 2.14fF
C2714 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<4> 0.01fF
C2715 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<14> 0.01fF
C2716 BU_3VX2_45|A vdd 0.06fF
C2717 raven_soc_0|flash_io1_oeb BU_3VX2_29|Q 0.01fF
C2718 raven_soc_0|flash_clk apllc03_1v8_0|CLK 0.01fF
C2719 BU_3VX2_47|Q vdd 2.70fF
C2720 vdd raven_padframe_0|VDDPADF_0|VDDR 0.71fF
C2721 markings_0|mask_copyright_0|m2_n208_960# markings_0|manufacturer_0|_alphabet_F_0|m2_0_0# 0.08fF
C2722 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<11> 1.25fF
C2723 raven_soc_0|gpio_out<0> VDD3V3 0.03fF
C2724 BU_3VX2_5|A BU_3VX2_6|Q 0.03fF
C2725 LS_3VX2_7|Q LS_3VX2_19|A 0.01fF
C2726 LS_3VX2_3|Q raven_soc_0|flash_io2_do 0.01fF
C2727 BU_3VX2_63|A raven_soc_0|flash_io0_do 0.01fF
C2728 LS_3VX2_14|Q LS_3VX2_22|A 0.31fF
C2729 VDD raven_padframe_0|FILLER50F_1|VDDR 0.71fF
C2730 BU_3VX2_28|A raven_soc_0|flash_io3_oeb 5.13fF
C2731 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<8> 0.42fF
C2732 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<12> 0.02fF
C2733 BU_3VX2_0|Q raven_soc_0|flash_io1_di 11.60fF
C2734 raven_soc_0|gpio_out<6> BU_3VX2_40|Q 0.01fF
C2735 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<15> 0.02fF
C2736 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<10> 0.01fF
C2737 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pullup<5> 0.05fF
C2738 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<7> 0.01fF
C2739 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<6> 0.01fF
C2740 raven_soc_0|gpio_out<9> raven_soc_0|ext_clk 0.01fF
C2741 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<13> 30.85fF
C2742 raven_soc_0|gpio_in<3> raven_soc_0|ext_clk 0.01fF
C2743 raven_soc_0|gpio_out<12> VDD3V3 0.07fF
C2744 raven_padframe_0|BBCUD4F_3|VDDR raven_padframe_0|BBCUD4F_3|GNDO 0.13fF
C2745 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<0> 0.01fF
C2746 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<19> 0.04fF
C2747 VDD raven_padframe_0|BBC4F_2|VDDR 0.71fF
C2748 BU_3VX2_7|A BU_3VX2_20|A 0.87fF
C2749 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<9> 0.01fF
C2750 BU_3VX2_2|A BU_3VX2_28|A 0.01fF
C2751 BU_3VX2_3|A BU_3VX2_3|Q 0.08fF
C2752 BU_3VX2_5|A raven_soc_0|flash_io2_di 0.03fF
C2753 LS_3VX2_12|A LS_3VX2_16|A 0.01fF
C2754 IN_3VX2_1|A raven_soc_0|gpio_pullup<14> 0.01fF
C2755 LOGIC0_3V_4|Q raven_soc_0|flash_io2_do 0.01fF
C2756 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<9> 0.87fF
C2757 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<13> 67.81fF
C2758 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<10> 121.55fF
C2759 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<8> 9.15fF
C2760 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pulldown<7> 0.02fF
C2761 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<14> 0.02fF
C2762 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pullup<13> 12.81fF
C2763 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<5> 0.01fF
C2764 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pulldown<6> 13.73fF
C2765 raven_soc_0|gpio_pullup<3> BU_3VX2_71|Q 0.01fF
C2766 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_15|PO 0.04fF
C2767 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_12|PO 0.04fF
C2768 raven_soc_0|gpio_pulldown<15> BU_3VX2_28|Q 0.01fF
C2769 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<18> 9.59fF
C2770 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<28> 0.01fF
C2771 BU_3VX2_6|Q BU_3VX2_68|Q 13.03fF
C2772 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<15> 0.39fF
C2773 BU_3VX2_16|Q BU_3VX2_5|Q 4.38fF
C2774 BU_3VX2_19|Q BU_3VX2_64|Q 0.01fF
C2775 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<8> 11.86fF
C2776 BU_3VX2_65|Q BU_3VX2_69|Q 4.81fF
C2777 BU_3VX2_68|Q BU_3VX2_7|Q 0.12fF
C2778 BU_3VX2_64|Q BU_3VX2_18|Q 0.02fF
C2779 BU_3VX2_5|Q BU_3VX2_30|Q 0.35fF
C2780 BU_3VX2_42|A BU_3VX2_42|Q 0.10fF
C2781 raven_padframe_0|FILLER20F_1|VDDO raven_padframe_0|FILLER20F_1|GNDO 2.28fF
C2782 BU_3VX2_10|A BU_3VX2_35|A 0.55fF
C2783 raven_padframe_0|BBC4F_2|VDDR LOGIC0_3V_4|Q 0.01fF
C2784 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<1> 7.10fF
C2785 BU_3VX2_18|A BU_3VX2_17|A 37.97fF
C2786 raven_spi_0|SDO LOGIC0_3V_2|Q 2.10fF
C2787 LS_3VX2_7|Q adc_low 0.12fF
C2788 raven_padframe_0|BBCUD4F_7|VDDO raven_padframe_0|BBCUD4F_7|GNDO 2.28fF
C2789 raven_padframe_0|CORNERESDF_1|VDDR raven_padframe_0|CORNERESDF_1|VDDO 0.06fF
C2790 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<12> 1.78fF
C2791 raven_soc_0|flash_io3_oeb BU_3VX2_33|Q 0.01fF
C2792 raven_soc_0|ram_addr<6> vdd 0.15fF
C2793 AMUX4_3V_1|SEL[0] BU_3VX2_54|Q 36.95fF
C2794 LOGIC0_3V_1|Q LOGIC0_3V_3|Q 7.38fF
C2795 VDD3V3 LS_3VX2_27|A 0.50fF
C2796 BU_3VX2_3|A BU_3VX2_22|A 2.79fF
C2797 BU_3VX2_35|A BU_3VX2_0|A 0.22fF
C2798 BU_3VX2_22|A BU_3VX2_15|A 2.48fF
C2799 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<6> 0.01fF
C2800 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<15> 0.01fF
C2801 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<11> 0.01fF
C2802 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<10> 0.01fF
C2803 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<9> 9.79fF
C2804 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<5> 0.02fF
C2805 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<12> 0.02fF
C2806 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<6> 2.42fF
C2807 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<7> 0.01fF
C2808 BU_3VX2_1|A VDD3V3 0.02fF
C2809 raven_soc_0|gpio_pulldown<2> BU_3VX2_40|Q 0.02fF
C2810 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<10> 1.17fF
C2811 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<31> 35.40fF
C2812 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<2> 11.57fF
C2813 raven_soc_0|ram_addr<9> raven_soc_0|ram_addr<3> 5.90fF
C2814 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<20> 0.01fF
C2815 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<29> 0.01fF
C2816 raven_soc_0|flash_io1_di raven_soc_0|flash_io3_di 132.18fF
C2817 BU_3VX2_13|Q BU_3VX2_36|Q 0.60fF
C2818 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<1> 0.72fF
C2819 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<13> 10.05fF
C2820 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<15> 8.00fF
C2821 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<17> 19.33fF
C2822 raven_soc_0|flash_io2_do raven_soc_0|flash_io1_oeb 44.88fF
C2823 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<22> 54.14fF
C2824 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<26> 0.01fF
C2825 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<25> 0.01fF
C2826 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<31> 11.38fF
C2827 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<19> 2.52fF
C2828 BU_3VX2_4|Q BU_3VX2_17|Q 2.42fF
C2829 BU_3VX2_46|A BU_3VX2_43|Q 0.02fF
C2830 raven_padframe_0|FILLER20F_5|VDDO raven_padframe_0|FILLER20F_5|GNDO 2.28fF
C2831 raven_spi_0|SDO raven_soc_0|flash_io0_do 0.50fF
C2832 BU_3VX2_38|A raven_soc_0|flash_io0_di 0.01fF
C2833 BU_3VX2_19|A raven_soc_0|flash_io3_do 0.01fF
C2834 raven_padframe_0|VDDPADF_1|VDDR vdd 0.71fF
C2835 LS_3VX2_10|Q VDD3V3 0.21fF
C2836 VDD raven_padframe_0|ICF_1|GNDO 0.07fF
C2837 BU_3VX2_63|Q BU_3VX2_35|Q 0.23fF
C2838 raven_soc_0|gpio_pulldown<13> BU_3VX2_29|Q 0.01fF
C2839 raven_soc_0|gpio_pullup<7> vdd 0.25fF
C2840 BU_3VX2_0|Q BU_3VX2_28|Q 0.02fF
C2841 raven_soc_0|gpio_outenb<0> BU_3VX2_26|Q 0.01fF
C2842 raven_soc_0|gpio_out<1> LOGIC0_3V_4|Q 0.01fF
C2843 LS_3VX2_12|Q LS_3VX2_5|Q 1.08fF
C2844 BU_3VX2_18|A BU_3VX2_12|A 3.07fF
C2845 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<3> 3.30fF
C2846 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<9> 0.01fF
C2847 raven_soc_0|gpio_pulldown<12> BU_3VX2_0|Q 0.01fF
C2848 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<10> 0.10fF
C2849 BU_3VX2_14|A raven_soc_0|flash_io3_oeb 0.01fF
C2850 raven_soc_0|gpio_pulldown<0> BU_3VX2_28|Q 0.01fF
C2851 raven_soc_0|gpio_outenb<2> BU_3VX2_27|Q 0.01fF
C2852 raven_soc_0|gpio_pullup<1> BU_3VX2_29|Q 0.01fF
C2853 raven_soc_0|gpio_pullup<5> VDD3V3 0.28fF
C2854 VDD3V3 BU_3VX2_54|A 0.05fF
C2855 raven_padframe_0|FILLER20FC_0|VDD3 raven_padframe_0|FILLER20FC_0|VDDR 0.71fF
C2856 LOGIC1_3V_2|Q LOGIC1_3V_0|Q 0.27fF
C2857 BU_3VX2_2|A BU_3VX2_14|A 1.08fF
C2858 BU_3VX2_38|A BU_3VX2_63|Q 0.02fF
C2859 BU_3VX2_0|A BU_3VX2_0|Q 0.09fF
C2860 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<12> 5.79fF
C2861 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<3> 19.16fF
C2862 BU_3VX2_31|A raven_soc_0|gpio_pullup<9> 0.01fF
C2863 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<7> 0.01fF
C2864 raven_padframe_0|BBCUD4F_14|VDDR raven_padframe_0|BBCUD4F_14|GNDO 0.13fF
C2865 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<20> 0.01fF
C2866 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<2> 7.76fF
C2867 raven_soc_0|gpio_pulldown<6> BU_3VX2_40|Q 0.57fF
C2868 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<14> 0.02fF
C2869 raven_soc_0|flash_io1_di raven_soc_0|irq_pin 0.01fF
C2870 BU_3VX2_16|Q BU_3VX2_28|Q 4.11fF
C2871 BU_3VX2_66|Q vdd 1.16fF
C2872 BU_3VX2_12|Q BU_3VX2_26|Q 0.03fF
C2873 BU_3VX2_6|Q BU_3VX2_24|Q 0.01fF
C2874 BU_3VX2_15|Q BU_3VX2_25|Q 3.54fF
C2875 BU_3VX2_73|Q LS_3VX2_15|A 0.01fF
C2876 LS_3VX2_22|A BU_3VX2_51|Q 7.86fF
C2877 BU_3VX2_30|Q BU_3VX2_28|Q 26.97fF
C2878 BU_3VX2_7|Q BU_3VX2_24|Q 0.02fF
C2879 BU_3VX2_64|Q BU_3VX2_27|Q 0.29fF
C2880 BU_3VX2_20|Q vdd 1.12fF
C2881 BU_3VX2_56|Q BU_3VX2_72|Q 1.09fF
C2882 BU_3VX2_65|Q BU_3VX2_29|Q 1.22fF
C2883 BU_3VX2_9|Q BU_3VX2_25|Q 1.11fF
C2884 LS_3VX2_17|A BU_3VX2_54|Q 8.64fF
C2885 BU_3VX2_33|Q apllc03_1v8_0|CLK 3.56fF
C2886 BU_3VX2_3|A BU_3VX2_21|A 1.14fF
C2887 BU_3VX2_21|A BU_3VX2_15|A 2.97fF
C2888 BU_3VX2_71|A BU_3VX2_17|A 0.01fF
C2889 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<5> 0.01fF
C2890 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<11> 0.01fF
C2891 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pullup<6> 7.97fF
C2892 raven_soc_0|ram_rdata<28> vdd 1.62fF
C2893 raven_soc_0|flash_io3_di BU_3VX2_28|Q 0.01fF
C2894 raven_soc_0|flash_io0_do BU_3VX2_26|Q 0.01fF
C2895 raven_soc_0|flash_io0_di BU_3VX2_23|Q 0.01fF
C2896 raven_soc_0|flash_io2_di BU_3VX2_24|Q 0.01fF
C2897 BU_3VX2_50|A vdd 0.06fF
C2898 raven_padframe_0|FILLER01F_1|GNDR raven_padframe_0|FILLER01F_1|VDDO 0.09fF
C2899 LOGIC0_3V_0|Q raven_soc_0|gpio_pulldown<15> 0.01fF
C2900 raven_padframe_0|FILLER50F_0|VDDR raven_padframe_0|FILLER50F_0|GNDR 0.68fF
C2901 raven_padframe_0|aregc01_3v3_1|VDDR raven_padframe_0|aregc01_3v3_1|GNDR 0.47fF
C2902 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<3> 2.52fF
C2903 LOGIC0_3V_1|Q VDD3V3 0.51fF
C2904 BU_3VX2_10|A raven_soc_0|flash_io3_di 0.04fF
C2905 BU_3VX2_8|A BU_3VX2_8|Q 0.08fF
C2906 LS_3VX2_14|A AMUX4_3V_1|SEL[0] 7.85fF
C2907 BU_3VX2_0|A BU_3VX2_30|Q 0.03fF
C2908 BU_3VX2_63|A raven_soc_0|flash_io1_di 0.01fF
C2909 LS_3VX2_7|Q LS_3VX2_22|A 0.01fF
C2910 IN_3VX2_1|A raven_soc_0|gpio_in<9> 0.01fF
C2911 LS_3VX2_4|Q LS_3VX2_19|A 0.01fF
C2912 raven_soc_0|gpio_outenb<11> BU_3VX2_40|Q 0.01fF
C2913 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pullup<5> 7.69fF
C2914 LS_3VX2_3|A raven_soc_0|flash_io3_oeb 0.01fF
C2915 raven_soc_0|gpio_outenb<10> raven_soc_0|ext_clk 0.01fF
C2916 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<11> 0.02fF
C2917 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<8> 0.01fF
C2918 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<7> 0.01fF
C2919 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<6> 0.01fF
C2920 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<13> 9.50fF
C2921 IN_3VX2_1|A BU_3VX2_42|Q 0.01fF
C2922 raven_soc_0|gpio_outenb<12> VDD3V3 0.07fF
C2923 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<11> 0.02fF
C2924 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<19> 2.88fF
C2925 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<0> 0.01fF
C2926 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<23> 0.07fF
C2927 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<20> 0.01fF
C2928 LS_3VX2_21|A adc0_data<5> 11.42fF
C2929 AMUX4_3V_3|AOUT AMUX4_3V_3|SEL[1] 0.36fF
C2930 VDD raven_padframe_0|ICF_2|GNDR 0.16fF
C2931 BU_3VX2_0|A raven_soc_0|flash_io3_di 9.53fF
C2932 BU_3VX2_35|A vdd 0.32fF
C2933 BU_3VX2_13|A raven_soc_0|flash_io2_di 0.01fF
C2934 raven_spi_0|sdo_enb raven_soc_0|flash_clk 0.42fF
C2935 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<13> 0.13fF
C2936 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<13> 29.53fF
C2937 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<9> 7.38fF
C2938 VDD raven_padframe_0|BBCUD4F_8|GNDR 0.16fF
C2939 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<14> 0.65fF
C2940 raven_soc_0|gpio_pulldown<5> BU_3VX2_71|Q 0.01fF
C2941 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<10> 18.74fF
C2942 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pulldown<6> 9.59fF
C2943 BU_3VX2_0|Q AMUX4_3V_4|SEL[0] 14.42fF
C2944 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<2> 0.01fF
C2945 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pulldown<7> 0.02fF
C2946 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<8> 4.69fF
C2947 raven_soc_0|gpio_pulldown<15> vdd 0.15fF
C2948 raven_soc_0|gpio_pulldown<14> BU_3VX2_26|Q 0.01fF
C2949 raven_soc_0|gpio_pulldown<11> BU_3VX2_24|Q 0.01fF
C2950 BU_3VX2_63|Q BU_3VX2_23|Q 0.01fF
C2951 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<12> 0.69fF
C2952 raven_soc_0|ram_wdata<1> raven_soc_0|ram_rdata<12> 2.86fF
C2953 VDD3V3 LS_3VX2_20|Q 0.18fF
C2954 BU_3VX2_8|A BU_3VX2_19|A 1.07fF
C2955 BU_3VX2_38|A BU_3VX2_5|A 1.60fF
C2956 BU_3VX2_71|A BU_3VX2_12|A 0.01fF
C2957 LS_3VX2_4|Q adc_low 0.12fF
C2958 raven_padframe_0|APR00DF_3|VDDR raven_padframe_0|APR00DF_3|VDDO 0.06fF
C2959 raven_soc_0|gpio_outenb<4> LS_3VX2_3|A 0.56fF
C2960 raven_soc_0|gpio_out<4> BU_3VX2_63|Q 0.01fF
C2961 raven_padframe_0|FILLER02F_1|GNDR raven_padframe_0|FILLER02F_1|VDDO 0.09fF
C2962 BU_3VX2_73|Q AMUX4_3V_1|SEL[1] 0.01fF
C2963 AMUX4_3V_1|SEL[0] BU_3VX2_56|Q 24.01fF
C2964 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<14> 0.01fF
C2965 BU_3VX2_35|A BU_3VX2_40|A 24.94fF
C2966 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<8> 0.01fF
C2967 LS_3VX2_8|A LS_3VX2_6|A 23.42fF
C2968 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<15> 0.01fF
C2969 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<10> 0.01fF
C2970 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<14> 3.68fF
C2971 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<11> 0.75fF
C2972 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<12> 0.51fF
C2973 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<12> 0.02fF
C2974 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<9> 6.23fF
C2975 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<5> 0.01fF
C2976 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<6> 0.01fF
C2977 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<7> 0.01fF
C2978 LS_3VX2_7|A BU_3VX2_73|Q 10.96fF
C2979 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<3> 9.41fF
C2980 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<31> 0.40fF
C2981 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<30> 20.39fF
C2982 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<9> 0.04fF
C2983 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<7> 9.71fF
C2984 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<20> 0.05fF
C2985 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<21> 0.01fF
C2986 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<24> 0.01fF
C2987 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<23> 0.01fF
C2988 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<18> 0.01fF
C2989 BU_3VX2_12|Q BU_3VX2_11|Q 67.20fF
C2990 BU_3VX2_66|Q BU_3VX2_70|Q 11.29fF
C2991 LS_3VX2_23|A BU_3VX2_7|Q 0.01fF
C2992 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<19> 22.57fF
C2993 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<25> 0.06fF
C2994 BU_3VX2_36|Q BU_3VX2_69|Q 2.02fF
C2995 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<27> 2.62fF
C2996 BU_3VX2_70|Q BU_3VX2_20|Q 0.01fF
C2997 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<2> 0.04fF
C2998 raven_soc_0|flash_io1_do raven_soc_0|flash_io3_oeb 121.64fF
C2999 BU_3VX2_3|Q BU_3VX2_17|Q 0.02fF
C3000 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<21> 0.02fF
C3001 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<13> 0.01fF
C3002 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<22> 0.01fF
C3003 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<14> 5.22fF
C3004 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<17> 0.01fF
C3005 BU_3VX2_32|Q BU_3VX2_67|Q 0.64fF
C3006 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<15> 6.21fF
C3007 BU_3VX2_72|Q BU_3VX2_29|Q 0.73fF
C3008 apllc03_1v8_0|CLK apllc03_1v8_0|B_CP 45.63fF
C3009 LOGIC0_3V_4|Q raven_soc_0|gpio_out<11> 0.01fF
C3010 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<13> 0.01fF
C3011 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<8> 0.01fF
C3012 AMUX4_3V_1|AIN1 AMUX4_3V_1|SEL[0] 0.02fF
C3013 BU_3VX2_2|A raven_soc_0|flash_io1_do 0.01fF
C3014 raven_spi_0|SDO raven_soc_0|flash_io1_di 1.43fF
C3015 VDD raven_padframe_0|BT4F_2|GNDR 0.16fF
C3016 LS_3VX2_14|A LS_3VX2_17|A 0.01fF
C3017 BU_3VX2_0|Q vdd 3.58fF
C3018 LS_3VX2_3|A apllc03_1v8_0|CLK 15.77fF
C3019 raven_soc_0|gpio_pulldown<10> BU_3VX2_26|Q 0.01fF
C3020 BU_3VX2_71|Q raven_soc_0|flash_io0_oeb 0.03fF
C3021 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<15> 15.21fF
C3022 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<16> 28.17fF
C3023 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<1> 17.82fF
C3024 BU_3VX2_10|A BU_3VX2_63|A 0.02fF
C3025 LS_3VX2_10|A BU_3VX2_59|Q 6.98fF
C3026 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<13> 0.47fF
C3027 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<15> 0.02fF
C3028 raven_soc_0|gpio_pulldown<0> vdd 0.32fF
C3029 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<11> 0.01fF
C3030 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<7> 4.99fF
C3031 raven_soc_0|gpio_out<2> BU_3VX2_23|Q 0.01fF
C3032 raven_soc_0|gpio_outenb<2> BU_3VX2_25|Q 0.91fF
C3033 BU_3VX2_63|A BU_3VX2_0|A 0.01fF
C3034 BU_3VX2_32|A BU_3VX2_33|A 1.54fF
C3035 BU_3VX2_40|A BU_3VX2_0|Q 2.09fF
C3036 LS_3VX2_14|Q LS_3VX2_5|A 0.18fF
C3037 IN_3VX2_1|A raven_soc_0|gpio_pullup<0> 0.01fF
C3038 IN_3VX2_1|A adc_high 0.28fF
C3039 LS_3VX2_6|A LS_3VX2_4|A 25.32fF
C3040 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<15> 0.67fF
C3041 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<5> 0.99fF
C3042 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<2> 1.92fF
C3043 BU_3VX2_31|A raven_soc_0|gpio_pulldown<9> 0.01fF
C3044 raven_soc_0|gpio_in<2> BU_3VX2_0|Q 0.01fF
C3045 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<9> 0.11fF
C3046 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<13> 16.79fF
C3047 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<5> 0.01fF
C3048 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<9> 0.01fF
C3049 BU_3VX2_24|A BU_3VX2_17|A 3.11fF
C3050 raven_soc_0|irq_pin comp_inp 25.15fF
C3051 BU_3VX2_16|Q vdd 0.71fF
C3052 BU_3VX2_35|Q BU_3VX2_24|Q 0.01fF
C3053 LS_3VX2_22|A BU_3VX2_49|Q 6.23fF
C3054 raven_soc_0|irq_pin BU_3VX2_44|Q 19.04fF
C3055 LS_3VX2_17|A BU_3VX2_56|Q 11.91fF
C3056 BU_3VX2_68|Q BU_3VX2_23|Q 2.87fF
C3057 BU_3VX2_30|Q vdd 1.61fF
C3058 BU_3VX2_5|Q BU_3VX2_26|Q 0.01fF
C3059 BU_3VX2_23|A IN_3VX2_1|A 5.44fF
C3060 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<7> 0.35fF
C3061 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_in<2> 6.23fF
C3062 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<17> 0.01fF
C3063 raven_soc_0|ram_wdata<21> raven_soc_0|ram_rdata<15> 0.93fF
C3064 raven_soc_0|ram_wdata<27> raven_soc_0|ram_rdata<1> 4.73fF
C3065 raven_soc_0|ram_wdata<22> raven_soc_0|ram_rdata<17> 0.04fF
C3066 raven_soc_0|ram_wdata<25> raven_soc_0|ram_addr<0> 0.01fF
C3067 raven_soc_0|flash_io3_di vdd 3.93fF
C3068 BU_3VX2_46|A LS_3VX2_27|Q 0.19fF
C3069 BU_3VX2_45|A LS_3VX2_21|Q 0.32fF
C3070 raven_soc_0|flash_io1_do apllc03_1v8_0|CLK 0.01fF
C3071 raven_soc_0|flash_io1_di BU_3VX2_26|Q 0.01fF
C3072 BU_3VX2_61|A BU_3VX2_60|Q 0.03fF
C3073 BU_3VX2_56|A BU_3VX2_59|Q 0.02fF
C3074 raven_soc_0|flash_io3_do BU_3VX2_27|Q 0.01fF
C3075 raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# raven_padframe_0|axtoc02_3v3_0|m4_55000_28769# 0.06fF
C3076 raven_padframe_0|axtoc02_3v3_0|m4_0_30133# raven_padframe_0|axtoc02_3v3_0|GNDR 0.15fF
C3077 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<7> 3.54fF
C3078 markings_0|date_0|_alphabet_1_1|m2_64_1376# markings_0|manufacturer_0|_alphabet_S_0|m2_32_224# 0.06fF
C3079 LS_3VX2_4|Q LS_3VX2_22|A 0.01fF
C3080 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<5> 0.85fF
C3081 raven_soc_0|gpio_pullup<11> BU_3VX2_40|Q 0.02fF
C3082 BU_3VX2_0|Q raven_soc_0|gpio_in<11> 0.33fF
C3083 raven_soc_0|gpio_pullup<12> VDD3V3 0.07fF
C3084 raven_soc_0|gpio_pullup<10> raven_soc_0|ext_clk 0.01fF
C3085 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<19> 31.38fF
C3086 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<0> 1.79fF
C3087 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<28> 24.27fF
C3088 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<20> 0.01fF
C3089 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<11> 5.86fF
C3090 BU_3VX2_36|Q BU_3VX2_29|Q 1.17fF
C3091 raven_soc_0|gpio_out<14> BU_3VX2_27|Q 0.01fF
C3092 BU_3VX2_71|Q BU_3VX2_29|Q 3.08fF
C3093 LS_3VX2_27|A adc0_data<5> 11.72fF
C3094 BU_3VX2_40|A raven_soc_0|flash_io3_di 0.39fF
C3095 BU_3VX2_18|A raven_soc_0|flash_clk 0.01fF
C3096 LOGIC0_3V_4|Q raven_soc_0|gpio_in<12> 0.08fF
C3097 BU_3VX2_31|A raven_soc_0|flash_io0_di 0.19fF
C3098 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<8> 5.31fF
C3099 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<6> 1.35fF
C3100 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<13> 0.57fF
C3101 raven_soc_0|gpio_in<2> raven_soc_0|flash_io3_di 0.22fF
C3102 BU_3VX2_0|Q raven_soc_0|gpio_outenb<9> 0.39fF
C3103 LS_3VX2_3|A raven_soc_0|gpio_outenb<8> 0.01fF
C3104 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<13> 6.17fF
C3105 BU_3VX2_33|A raven_soc_0|flash_io2_oeb 0.01fF
C3106 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pulldown<6> 0.02fF
C3107 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<14> 0.02fF
C3108 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<16> 1.86fF
C3109 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<2> 60.29fF
C3110 BU_3VX2_0|Q BU_3VX2_70|Q 0.01fF
C3111 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<8> 4.60fF
C3112 AMUX2_3V_0|SEL BU_3VX2_50|Q 6.21fF
C3113 LS_3VX2_13|A AMUX4_3V_4|AIN2 0.63fF
C3114 raven_padframe_0|BBCUD4F_0|VDDR raven_padframe_0|BBCUD4F_0|VDDO 0.06fF
C3115 BU_3VX2_24|A BU_3VX2_12|A 1.73fF
C3116 BU_3VX2_9|A BU_3VX2_18|A 1.36fF
C3117 BU_3VX2_38|A BU_3VX2_13|A 1.02fF
C3118 BU_3VX2_5|A BU_3VX2_4|Q 0.16fF
C3119 raven_padframe_0|ICFC_0|VDDR raven_padframe_0|ICFC_0|VDDO 0.06fF
C3120 LOGIC0_3V_4|Q raven_padframe_0|ICFC_2|PO 0.04fF
C3121 raven_soc_0|irq_pin vdd 5.66fF
C3122 AMUX4_3V_3|SEL[0] comp_inp 0.02fF
C3123 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<15> 0.01fF
C3124 BU_3VX2_16|A BU_3VX2_17|A 39.99fF
C3125 LS_3VX2_10|A AMUX2_3V_0|SEL 11.06fF
C3126 BU_3VX2_17|A BU_3VX2_29|A 1.77fF
C3127 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_out<3> 2.69fF
C3128 BU_3VX2_26|A LOGIC0_3V_2|Q 0.01fF
C3129 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<6> 0.03fF
C3130 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<7> 0.02fF
C3131 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<10> 27.59fF
C3132 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<5> 0.68fF
C3133 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<4> 0.55fF
C3134 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<11> 9.88fF
C3135 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<6> 0.01fF
C3136 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<14> 0.02fF
C3137 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<11> 6.36fF
C3138 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<12> 0.02fF
C3139 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<2> 0.01fF
C3140 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<26> 4.02fF
C3141 raven_soc_0|flash_io3_do raven_soc_0|flash_io2_oeb 49.20fF
C3142 BU_3VX2_15|Q BU_3VX2_37|Q 15.19fF
C3143 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<30> 4.69fF
C3144 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<23> 13.31fF
C3145 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<10> 0.11fF
C3146 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<21> 17.98fF
C3147 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<14> 4.41fF
C3148 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<7> 0.64fF
C3149 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<2> 0.72fF
C3150 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<12> 1.34fF
C3151 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<9> 0.10fF
C3152 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<17> 0.02fF
C3153 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<0> 0.01fF
C3154 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<4> 40.04fF
C3155 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<25> 5.65fF
C3156 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<7> 10.90fF
C3157 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<14> 0.02fF
C3158 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<10> 0.01fF
C3159 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<4> 0.01fF
C3160 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<15> 0.01fF
C3161 BU_3VX2_32|Q BU_3VX2_65|Q 24.03fF
C3162 BU_3VX2_11|Q BU_3VX2_5|Q 8.38fF
C3163 BU_3VX2_14|Q BU_3VX2_22|Q 4.98fF
C3164 BU_3VX2_70|Q BU_3VX2_30|Q 2.41fF
C3165 AMUX4_3V_4|SEL[0] AMUX4_3V_3|SEL[0] 168.51fF
C3166 BU_3VX2_37|Q BU_3VX2_9|Q 4.49fF
C3167 BU_3VX2_26|Q BU_3VX2_28|Q 93.44fF
C3168 BU_3VX2_24|Q BU_3VX2_23|Q 359.66fF
C3169 BU_3VX2_25|Q apllc03_1v8_0|B_VCO 0.83fF
C3170 BU_3VX2_23|A BU_3VX2_25|A 19.83fF
C3171 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<15> 0.01fF
C3172 raven_padframe_0|CORNERESDF_0|VDDR raven_padframe_0|CORNERESDF_0|VDDO 0.06fF
C3173 BU_3VX2_11|A LOGIC0_3V_2|Q 0.01fF
C3174 LOGIC0_3V_3|Q LOGIC0_3V_2|Q 22.13fF
C3175 raven_padframe_0|aregc01_3v3_0|VDDO raven_padframe_0|aregc01_3v3_0|GNDO 1.69fF
C3176 BU_3VX2_6|A raven_soc_0|flash_io3_do 0.02fF
C3177 BU_3VX2_63|A vdd 0.09fF
C3178 BU_3VX2_64|A BU_3VX2_64|Q 0.08fF
C3179 raven_soc_0|gpio_in<2> raven_soc_0|irq_pin 0.13fF
C3180 raven_soc_0|gpio_pulldown<12> BU_3VX2_26|Q 0.01fF
C3181 raven_soc_0|ser_rx AMUX4_3V_4|AIN2 11.75fF
C3182 BU_3VX2_71|Q raven_soc_0|flash_io2_do 0.01fF
C3183 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<1> 27.28fF
C3184 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<13> 6.64fF
C3185 raven_soc_0|ser_tx BU_3VX2_59|Q 8.51fF
C3186 raven_soc_0|ram_rdata<31> apllc03_1v8_0|CLK 3.51fF
C3187 LS_3VX2_10|A BU_3VX2_61|Q 0.01fF
C3188 BU_3VX2_11|A BU_3VX2_12|Q 0.03fF
C3189 LS_3VX2_24|A BU_3VX2_59|Q 0.02fF
C3190 BU_3VX2_69|A BU_3VX2_66|Q 0.02fF
C3191 BU_3VX2_26|A raven_soc_0|flash_io0_do 2.66fF
C3192 LS_3VX2_6|A vdd 3.64fF
C3193 VDD raven_padframe_0|aregc01_3v3_1|GNDR 0.10fF
C3194 raven_soc_0|gpio_pulldown<8> BU_3VX2_40|Q 0.21fF
C3195 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<8> 0.01fF
C3196 BU_3VX2_0|Q raven_soc_0|ram_rdata<24> 0.02fF
C3197 raven_soc_0|gpio_pulldown<1> BU_3VX2_27|Q 0.01fF
C3198 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<6> 0.01fF
C3199 BU_3VX2_63|A BU_3VX2_40|A 0.13fF
C3200 BU_3VX2_16|A BU_3VX2_12|A 4.98fF
C3201 BU_3VX2_18|A BU_3VX2_28|A 2.14fF
C3202 BU_3VX2_29|A BU_3VX2_12|A 0.01fF
C3203 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<3> 0.69fF
C3204 AMUX4_3V_3|AOUT raven_soc_0|flash_io1_oeb 2.52fF
C3205 BU_3VX2_22|A raven_soc_0|flash_io0_di 0.01fF
C3206 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<9> 0.01fF
C3207 BU_3VX2_71|A raven_soc_0|flash_clk 0.01fF
C3208 raven_soc_0|gpio_in<3> raven_soc_0|flash_io2_di 2.66fF
C3209 BU_3VX2_63|Q raven_soc_0|gpio_out<8> 0.41fF
C3210 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<13> 34.10fF
C3211 BU_3VX2_11|A raven_soc_0|flash_io0_do 0.01fF
C3212 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<10> 8.82fF
C3213 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<3> 4.24fF
C3214 raven_soc_0|flash_csb raven_soc_0|flash_io3_oeb 40.85fF
C3215 LOGIC0_3V_0|Q raven_spi_0|SDO 3.66fF
C3216 raven_soc_0|gpio_in<11> raven_soc_0|irq_pin 0.03fF
C3217 AMUX4_3V_3|SEL[0] vdd 2.80fF
C3218 VDD raven_padframe_0|BBCUD4F_11|VDDR 0.71fF
C3219 BU_3VX2_9|A BU_3VX2_71|A 0.02fF
C3220 BU_3VX2_37|A BU_3VX2_12|A 1.30fF
C3221 LS_3VX2_3|Q BU_3VX2_17|A 0.01fF
C3222 BU_3VX2_5|A BU_3VX2_31|A 0.01fF
C3223 raven_soc_0|gpio_pullup<2> BU_3VX2_0|Q 0.01fF
C3224 BU_3VX2_2|A raven_soc_0|flash_csb 0.01fF
C3225 BU_3VX2_31|A raven_soc_0|gpio_out<2> 0.01fF
C3226 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<0> 9.16fF
C3227 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<17> 6.94fF
C3228 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<1> 0.06fF
C3229 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<15> 1.83fF
C3230 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<25> 0.01fF
C3231 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<27> 0.01fF
C3232 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<31> 0.01fF
C3233 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<22> 0.01fF
C3234 raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<29> 27.55fF
C3235 raven_soc_0|ram_wdata<17> raven_soc_0|ram_rdata<13> 0.02fF
C3236 raven_soc_0|ram_wdata<26> raven_soc_0|ram_rdata<1> 2.74fF
C3237 raven_soc_0|ram_wdata<14> raven_soc_0|ram_rdata<15> 0.07fF
C3238 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<31> 6.55fF
C3239 AMUX4_3V_0|SEL[1] BU_3VX2_45|Q 35.77fF
C3240 raven_soc_0|gpio_in<10> apllc03_1v8_0|CLK 0.02fF
C3241 BU_3VX2_50|A LS_3VX2_21|Q 0.12fF
C3242 BU_3VX2_51|A BU_3VX2_42|A 0.12fF
C3243 BU_3VX2_48|A BU_3VX2_44|A 0.59fF
C3244 BU_3VX2_49|A BU_3VX2_43|A 0.32fF
C3245 BU_3VX2_61|A BU_3VX2_62|Q 0.14fF
C3246 raven_soc_0|gpio_out<15> BU_3VX2_23|Q 0.01fF
C3247 raven_soc_0|flash_io3_do BU_3VX2_25|Q 0.01fF
C3248 BU_3VX2_45|Q BU_3VX2_51|Q 16.76fF
C3249 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<3> 3.52fF
C3250 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<0> 4.97fF
C3251 raven_padframe_0|BBCUD4F_11|VDDR LOGIC0_3V_4|Q 0.01fF
C3252 BU_3VX2_25|A IN_3VX2_1|A 6.88fF
C3253 LS_3VX2_10|Q LS_3VX2_24|Q 0.01fF
C3254 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_in<0> 0.01fF
C3255 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<2> 0.52fF
C3256 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<5> 0.28fF
C3257 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<11> 0.01fF
C3258 raven_padframe_0|axtoc02_3v3_0|m4_55000_31172# raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# 0.03fF
C3259 raven_padframe_0|axtoc02_3v3_0|m4_0_29333# raven_padframe_0|axtoc02_3v3_0|m4_0_22024# 0.02fF
C3260 BU_3VX2_63|Q raven_soc_0|gpio_out<6> 0.01fF
C3261 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<14> 18.82fF
C3262 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<5> 0.01fF
C3263 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<9> 4.25fF
C3264 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<7> 4.63fF
C3265 markings_0|date_0|_alphabet_1_1|m2_64_1376# markings_0|date_0|_alphabet_0_0|m2_0_208# 0.61fF
C3266 raven_soc_0|gpio_out<1> BU_3VX2_71|Q 0.01fF
C3267 LS_3VX2_14|A BU_3VX2_42|Q 7.94fF
C3268 BU_3VX2_66|A BU_3VX2_64|Q 0.03fF
C3269 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<12> 17.31fF
C3270 LS_3VX2_3|A raven_soc_0|gpio_in<15> 0.01fF
C3271 adc_high BU_3VX2_54|Q 0.17fF
C3272 raven_soc_0|gpio_outenb<0> VDD3V3 0.03fF
C3273 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<9> 0.02fF
C3274 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<8> 3.93fF
C3275 raven_soc_0|gpio_pulldown<4> raven_soc_0|ext_clk 0.01fF
C3276 raven_soc_0|gpio_pullup<14> BU_3VX2_29|Q 0.01fF
C3277 raven_soc_0|gpio_outenb<13> BU_3VX2_28|Q 0.01fF
C3278 raven_soc_0|gpio_out<14> BU_3VX2_25|Q 0.01fF
C3279 BU_3VX2_11|Q BU_3VX2_28|Q 6.44fF
C3280 BU_3VX2_4|Q BU_3VX2_24|Q 7.60fF
C3281 BU_3VX2_10|A BU_3VX2_11|Q 0.03fF
C3282 BU_3VX2_8|A raven_soc_0|flash_io2_oeb 0.01fF
C3283 BU_3VX2_20|A raven_soc_0|flash_io3_oeb 0.01fF
C3284 LS_3VX2_11|Q VDD3V3 0.21fF
C3285 raven_padframe_0|BBC4F_2|VDDR raven_padframe_0|BBC4F_2|GNDO 0.13fF
C3286 VDD raven_padframe_0|ICF_0|GNDR 0.16fF
C3287 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pulldown<6> 0.97fF
C3288 raven_spi_0|sdo_enb raven_soc_0|flash_io1_do 0.71fF
C3289 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<13> 0.02fF
C3290 BU_3VX2_27|A raven_soc_0|flash_io3_do 0.01fF
C3291 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<13> 40.79fF
C3292 LOGIC0_3V_2|Q VDD3V3 0.28fF
C3293 AMUX2_3V_0|SEL BU_3VX2_48|Q 5.15fF
C3294 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<23> 24.29fF
C3295 BU_3VX2_41|A BU_3VX2_46|A 7.98fF
C3296 BU_3VX2_8|A BU_3VX2_6|A 8.03fF
C3297 BU_3VX2_73|A analog_out 0.02fF
C3298 LS_3VX2_3|Q BU_3VX2_12|A 0.01fF
C3299 BU_3VX2_21|A raven_soc_0|flash_io0_di 0.15fF
C3300 LS_3VX2_12|A LS_3VX2_19|A 0.01fF
C3301 BU_3VX2_5|A BU_3VX2_3|Q 0.03fF
C3302 raven_soc_0|gpio_out<0> BU_3VX2_27|Q 0.07fF
C3303 LS_3VX2_12|A BU_3VX2_52|Q 8.28fF
C3304 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<7> 0.01fF
C3305 BU_3VX2_17|A raven_soc_0|flash_io1_oeb 0.01fF
C3306 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<8> 1.16fF
C3307 AMUX2_3V_0|SEL raven_soc_0|ser_tx 0.01fF
C3308 raven_soc_0|gpio_in<0> apllc03_1v8_0|CLK 0.03fF
C3309 raven_soc_0|flash_csb apllc03_1v8_0|CLK 0.01fF
C3310 raven_soc_0|gpio_out<12> BU_3VX2_27|Q 0.01fF
C3311 BU_3VX2_57|A BU_3VX2_56|Q 0.03fF
C3312 BU_3VX2_52|A BU_3VX2_55|Q 0.02fF
C3313 raven_soc_0|gpio_in<7> raven_padframe_0|BBCUD4F_7|PO 0.04fF
C3314 BU_3VX2_7|A BU_3VX2_35|A 0.84fF
C3315 BU_3VX2_23|A BU_3VX2_4|A 0.01fF
C3316 LS_3VX2_6|Q LS_3VX2_10|Q 10.89fF
C3317 BU_3VX2_18|A BU_3VX2_14|A 5.53fF
C3318 BU_3VX2_71|A BU_3VX2_28|A 0.01fF
C3319 BU_3VX2_0|A BU_3VX2_36|A 8.82fF
C3320 LS_3VX2_24|A AMUX2_3V_0|SEL 61.24fF
C3321 BU_3VX2_64|A BU_3VX2_33|A 2.57fF
C3322 raven_soc_0|gpio_pulldown<2> BU_3VX2_63|Q 0.01fF
C3323 BU_3VX2_69|A BU_3VX2_0|Q 1.21fF
C3324 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<6> 0.19fF
C3325 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<12> 1.73fF
C3326 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<11> 8.94fF
C3327 LS_3VX2_3|A raven_soc_0|gpio_out<13> 0.01fF
C3328 BU_3VX2_0|Q raven_soc_0|gpio_outenb<14> 0.01fF
C3329 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<5> 0.01fF
C3330 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<15> 0.02fF
C3331 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<11> 8.50fF
C3332 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<5> 0.01fF
C3333 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<25> 0.28fF
C3334 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<8> 0.26fF
C3335 AMUX4_3V_3|SEL[1] BU_3VX2_10|Q 0.09fF
C3336 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<7> 3.12fF
C3337 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<14> 0.44fF
C3338 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<18> 0.27fF
C3339 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<12> 0.03fF
C3340 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<8> 0.15fF
C3341 AMUX4_3V_3|SEL[1] BU_3VX2_2|Q 6.75fF
C3342 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<1> 0.01fF
C3343 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<2> 0.21fF
C3344 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<4> 0.02fF
C3345 raven_soc_0|ext_clk raven_soc_0|flash_io2_di 56.48fF
C3346 BU_3VX2_3|Q BU_3VX2_68|Q 5.62fF
C3347 BU_3VX2_14|Q BU_3VX2_31|Q 0.02fF
C3348 raven_soc_0|flash_io0_do VDD3V3 12.14fF
C3349 vdd BU_3VX2_26|Q 2.19fF
C3350 BU_3VX2_22|A BU_3VX2_5|A 0.92fF
C3351 LS_3VX2_8|Q LS_3VX2_10|Q 1.24fF
C3352 raven_padframe_0|aregc01_3v3_0|m4_92500_29057# raven_padframe_0|aregc01_3v3_0|VDDO 0.04fF
C3353 raven_padframe_0|aregc01_3v3_0|m4_92500_29333# raven_padframe_0|aregc01_3v3_0|GNDO 0.12fF
C3354 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<6> 0.28fF
C3355 AMUX4_3V_1|AIN1 BU_3VX2_57|A 0.02fF
C3356 LS_3VX2_7|A BU_3VX2_43|Q 0.10fF
C3357 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<21> 0.02fF
C3358 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<10> 3.62fF
C3359 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<20> 0.01fF
C3360 raven_soc_0|ser_tx BU_3VX2_61|Q 11.62fF
C3361 raven_soc_0|ram_rdata<10> vdd 0.15fF
C3362 raven_soc_0|ram_rdata<30> apllc03_1v8_0|CLK 3.23fF
C3363 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<3> 2.62fF
C3364 BU_3VX2_15|A BU_3VX2_15|Q 0.08fF
C3365 LS_3VX2_10|A LS_3VX2_15|A 0.02fF
C3366 AMUX4_3V_0|AIN1 LS_3VX2_20|Q 0.96fF
C3367 BU_3VX2_12|A raven_soc_0|flash_io1_oeb 0.01fF
C3368 LS_3VX2_24|A BU_3VX2_61|Q 0.02fF
C3369 BU_3VX2_31|A BU_3VX2_24|Q 25.75fF
C3370 BU_3VX2_26|A raven_soc_0|flash_io1_di 0.01fF
C3371 BU_3VX2_0|Q LS_3VX2_2|A 6.01fF
C3372 raven_soc_0|gpio_pulldown<1> BU_3VX2_25|Q 0.01fF
C3373 raven_soc_0|gpio_pulldown<11> raven_soc_0|ext_clk 0.01fF
C3374 IN_3VX2_1|A BU_3VX2_54|Q 0.01fF
C3375 raven_soc_0|gpio_pulldown<14> VDD3V3 0.07fF
C3376 raven_soc_0|gpio_in<2> BU_3VX2_26|Q 0.01fF
C3377 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<10> 9.05fF
C3378 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<31> 0.61fF
C3379 BU_3VX2_32|Q BU_3VX2_36|Q 3.21fF
C3380 raven_padframe_0|FILLER10F_1|VDDR raven_padframe_0|FILLER10F_1|GNDO 0.13fF
C3381 BU_3VX2_32|A BU_3VX2_1|A 6.92fF
C3382 BU_3VX2_24|A raven_soc_0|flash_clk 4.03fF
C3383 LS_3VX2_4|Q LS_3VX2_5|A 0.16fF
C3384 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<5> 0.17fF
C3385 raven_soc_0|gpio_out<0> raven_soc_0|flash_io2_oeb 0.93fF
C3386 BU_3VX2_11|A raven_soc_0|flash_io1_di 0.01fF
C3387 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<6> 0.01fF
C3388 LOGIC0_3V_1|Q LOGIC1_3V_3|Q 0.14fF
C3389 BU_3VX2_24|A BU_3VX2_9|A 0.01fF
C3390 BU_3VX2_8|A BU_3VX2_27|A 0.01fF
C3391 BU_3VX2_4|A IN_3VX2_1|A 0.01fF
C3392 BU_3VX2_66|A BU_3VX2_33|A 1.65fF
C3393 BU_3VX2_31|A BU_3VX2_13|A 0.01fF
C3394 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_out<2> 19.82fF
C3395 LS_3VX2_12|A BU_3VX2_58|Q 0.01fF
C3396 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<8> 0.01fF
C3397 raven_soc_0|gpio_out<11> BU_3VX2_71|Q 0.01fF
C3398 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<8> 3.74fF
C3399 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<9> 0.01fF
C3400 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<6> 10.11fF
C3401 raven_soc_0|ram_wdata<1> raven_soc_0|ram_rdata<16> 1.31fF
C3402 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<31> 202.25fF
C3403 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<22> 0.01fF
C3404 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<1> 4.14fF
C3405 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<17> 0.01fF
C3406 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<19> 0.01fF
C3407 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<13> 0.01fF
C3408 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<29> 0.01fF
C3409 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<26> 0.01fF
C3410 raven_soc_0|gpio_in<9> BU_3VX2_29|Q 0.01fF
C3411 raven_soc_0|gpio_in<13> apllc03_1v8_0|CLK 0.02fF
C3412 LS_3VX2_15|Q LS_3VX2_16|A 0.19fF
C3413 AMUX4_3V_1|SEL[0] AMUX4_3V_4|AIN2 0.01fF
C3414 raven_soc_0|gpio_in<11> BU_3VX2_26|Q 0.01fF
C3415 AMUX4_3V_0|SEL[0] BU_3VX2_44|Q 34.01fF
C3416 raven_soc_0|gpio_in<8> BU_3VX2_28|Q 0.01fF
C3417 BU_3VX2_45|Q BU_3VX2_49|Q 25.07fF
C3418 BU_3VX2_21|A BU_3VX2_5|A 1.25fF
C3419 LS_3VX2_22|Q aopac01_3v3_0|IB 0.10fF
C3420 BU_3VX2_71|A BU_3VX2_14|A 0.01fF
C3421 raven_padframe_0|aregc01_3v3_1|m4_0_28769# raven_padframe_0|aregc01_3v3_1|m4_0_22024# 0.03fF
C3422 raven_padframe_0|aregc01_3v3_1|m4_92500_30133# raven_padframe_0|aregc01_3v3_1|m4_92500_29057# 0.01fF
C3423 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<7> 0.01fF
C3424 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<15> 340.91fF
C3425 BU_3VX2_63|Q raven_soc_0|gpio_outenb<11> 0.01fF
C3426 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<10> 10.70fF
C3427 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<6> 0.01fF
C3428 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<9> 9.76fF
C3429 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<14> 0.16fF
C3430 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<6> 0.11fF
C3431 LS_3VX2_7|A BU_3VX2_50|Q 0.11fF
C3432 LS_3VX2_3|A raven_soc_0|gpio_in<14> 0.01fF
C3433 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<8> 0.01fF
C3434 raven_soc_0|gpio_pulldown<10> VDD3V3 0.07fF
C3435 adc_high BU_3VX2_56|Q 0.11fF
C3436 raven_soc_0|gpio_outenb<13> vdd 0.21fF
C3437 raven_soc_0|gpio_outenb<9> BU_3VX2_26|Q 0.01fF
C3438 raven_soc_0|gpio_pullup<13> BU_3VX2_28|Q 0.01fF
C3439 raven_soc_0|gpio_out<10> BU_3VX2_23|Q 0.01fF
C3440 BU_3VX2_70|Q BU_3VX2_26|Q 0.31fF
C3441 BU_3VX2_11|Q vdd 1.19fF
C3442 raven_soc_0|flash_io2_di raven_padframe_0|BBC4F_3|PO 0.04fF
C3443 BU_3VX2_3|Q BU_3VX2_24|Q 0.01fF
C3444 BU_3VX2_14|Q apllc03_1v8_0|CLK 0.01fF
C3445 BU_3VX2_7|A raven_soc_0|flash_io3_di 0.01fF
C3446 LS_3VX2_10|A AMUX4_3V_1|SEL[1] 23.63fF
C3447 raven_padframe_0|BT4F_2|VDDR raven_padframe_0|BT4F_2|VDDO 0.06fF
C3448 BU_3VX2_18|A raven_soc_0|flash_io1_do 0.01fF
C3449 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<10> 0.57fF
C3450 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<7> 2.20fF
C3451 BU_3VX2_31|A raven_soc_0|gpio_out<15> 0.01fF
C3452 analog_out comp_inp 9.44fF
C3453 raven_soc_0|gpio_outenb<2> BU_3VX2_40|Q 1.80fF
C3454 LS_3VX2_3|A raven_soc_0|gpio_pullup<6> 0.17fF
C3455 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<13> 19.32fF
C3456 BU_3VX2_0|Q raven_soc_0|ram_wdata<27> 0.02fF
C3457 BU_3VX2_36|A vdd 0.79fF
C3458 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<20> 4.73fF
C3459 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<0> 0.33fF
C3460 BU_3VX2_47|A adc0_data<5> 0.15fF
C3461 raven_padframe_0|APR00DF_6|VDDR raven_padframe_0|APR00DF_6|GNDO 0.13fF
C3462 raven_padframe_0|APR00DF_6|GNDR raven_padframe_0|APR00DF_6|VDDO 0.09fF
C3463 raven_padframe_0|BBCUD4F_11|GNDR raven_padframe_0|BBCUD4F_11|VDDO 0.09fF
C3464 raven_padframe_0|APR00DF_4|GNDR raven_padframe_0|APR00DF_4|GNDO 0.81fF
C3465 LS_3VX2_10|A LS_3VX2_7|A 32.36fF
C3466 BU_3VX2_10|A BU_3VX2_26|A 0.01fF
C3467 AMUX4_3V_1|AIN1 adc_high 0.22fF
C3468 BU_3VX2_23|A raven_soc_0|flash_io0_oeb 3.38fF
C3469 LS_3VX2_12|A LS_3VX2_22|A 18.27fF
C3470 BU_3VX2_37|A BU_3VX2_2|Q 0.03fF
C3471 BU_3VX2_16|A raven_soc_0|flash_clk 0.01fF
C3472 raven_soc_0|gpio_out<0> BU_3VX2_25|Q 0.01fF
C3473 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<13> 0.01fF
C3474 BU_3VX2_29|A raven_soc_0|flash_clk 12.80fF
C3475 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<7> 0.01fF
C3476 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<6> 0.01fF
C3477 VDD raven_padframe_0|APR00DF_4|GNDO 0.07fF
C3478 raven_soc_0|gpio_out<12> BU_3VX2_25|Q 0.01fF
C3479 raven_soc_0|gpio_outenb<12> BU_3VX2_27|Q 0.01fF
C3480 BU_3VX2_73|Q LS_3VX2_20|A 18.70fF
C3481 raven_soc_0|ext_clk BU_3VX2_57|Q 0.01fF
C3482 BU_3VX2_24|A BU_3VX2_28|A 9.71fF
C3483 VDD3V3 raven_padframe_0|VDDORPADF_2|GNDR 0.78fF
C3484 BU_3VX2_9|A BU_3VX2_16|A 1.78fF
C3485 BU_3VX2_10|A BU_3VX2_11|A 22.43fF
C3486 BU_3VX2_9|A BU_3VX2_29|A 0.01fF
C3487 BU_3VX2_0|A BU_3VX2_26|A 0.01fF
C3488 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<1> 2.44fF
C3489 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<3> 5.21fF
C3490 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<9> 0.83fF
C3491 BU_3VX2_37|A raven_soc_0|flash_clk 0.01fF
C3492 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<6> 0.01fF
C3493 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<8> 0.36fF
C3494 LS_3VX2_3|A raven_soc_0|gpio_outenb<15> 0.01fF
C3495 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<5> 0.01fF
C3496 BU_3VX2_0|Q raven_soc_0|gpio_pullup<15> 0.01fF
C3497 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<11> 6.39fF
C3498 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<10> 0.19fF
C3499 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<14> 0.39fF
C3500 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<9> 0.02fF
C3501 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<10> 7.78fF
C3502 raven_soc_0|gpio_in<15> raven_soc_0|gpio_in<10> 10.15fF
C3503 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<1> 1.05fF
C3504 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<0> 1.88fF
C3505 AMUX4_3V_3|SEL[1] BU_3VX2_33|Q 1.07fF
C3506 raven_soc_0|flash_io1_di VDD3V3 9.22fF
C3507 AMUX4_3V_0|SEL[0] vdd 3.26fF
C3508 AMUX4_3V_4|AIN2 LS_3VX2_17|A 0.01fF
C3509 BU_3VX2_9|A BU_3VX2_37|A 0.94fF
C3510 raven_padframe_0|POWERCUTVDD3FC_0|VDDR LOGIC0_3V_4|Q 0.01fF
C3511 BU_3VX2_22|A BU_3VX2_13|A 1.77fF
C3512 BU_3VX2_25|A BU_3VX2_4|A 0.01fF
C3513 BU_3VX2_0|A BU_3VX2_11|A 0.01fF
C3514 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<4> 0.01fF
C3515 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<11> 0.50fF
C3516 raven_padframe_0|aregc01_3v3_0|m4_92500_29333# raven_padframe_0|aregc01_3v3_0|m4_92500_29057# 0.11fF
C3517 raven_padframe_0|aregc01_3v3_0|m4_92500_30133# raven_padframe_0|aregc01_3v3_0|m4_92500_28769# 0.01fF
C3518 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<7> 0.71fF
C3519 BU_3VX2_38|A raven_soc_0|ext_clk 0.01fF
C3520 BU_3VX2_73|A VDD3V3 0.10fF
C3521 BU_3VX2_68|A BU_3VX2_69|Q 0.03fF
C3522 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<28> 11.24fF
C3523 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<7> 0.98fF
C3524 BU_3VX2_71|Q raven_soc_0|gpio_in<12> 0.02fF
C3525 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<2> 0.03fF
C3526 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<11> 9.64fF
C3527 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<15> 0.11fF
C3528 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<17> 0.02fF
C3529 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<26> 0.01fF
C3530 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<19> 0.02fF
C3531 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<13> 0.02fF
C3532 raven_soc_0|gpio_out<8> raven_soc_0|gpio_out<15> 0.02fF
C3533 raven_soc_0|ram_addr<3> vdd 0.22fF
C3534 raven_soc_0|ser_tx LS_3VX2_15|A 14.59fF
C3535 AMUX4_3V_0|SEL[1] LS_3VX2_21|A 6.99fF
C3536 LS_3VX2_21|A BU_3VX2_51|Q 33.98fF
C3537 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<15> 0.01fF
C3538 IN_3VX2_1|Q BU_3VX2_43|Q 1.54fF
C3539 LS_3VX2_8|A VDD3V3 0.52fF
C3540 VDD raven_padframe_0|BBC4F_1|GNDO 0.07fF
C3541 LS_3VX2_24|A LS_3VX2_15|A 0.02fF
C3542 raven_soc_0|gpio_pullup<0> BU_3VX2_29|Q 0.01fF
C3543 IN_3VX2_1|A BU_3VX2_56|Q 0.01fF
C3544 raven_soc_0|gpio_pulldown<2> BU_3VX2_24|Q 0.01fF
C3545 raven_soc_0|gpio_outenb<1> apllc03_1v8_0|CLK 0.01fF
C3546 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_outenb<13> 1.54fF
C3547 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<5> 0.04fF
C3548 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<10> 0.13fF
C3549 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<7> 0.23fF
C3550 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<31> 0.03fF
C3551 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<24> 161.63fF
C3552 BU_3VX2_70|Q BU_3VX2_11|Q 0.60fF
C3553 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<6> 0.46fF
C3554 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<9> 0.07fF
C3555 raven_soc_0|ram_wdata<20> raven_soc_0|ram_addr<2> 0.01fF
C3556 BU_3VX2_7|A BU_3VX2_63|A 0.01fF
C3557 BU_3VX2_71|A raven_soc_0|flash_io1_do 0.01fF
C3558 raven_soc_0|gpio_pullup<2> BU_3VX2_26|Q 0.01fF
C3559 LS_3VX2_3|Q raven_soc_0|flash_clk 0.01fF
C3560 BU_3VX2_67|A BU_3VX2_67|Q 0.08fF
C3561 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<15> 9.16fF
C3562 VDD raven_padframe_0|FILLER20F_0|GNDR 0.16fF
C3563 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<3> 1.95fF
C3564 IN_3VX2_1|A raven_soc_0|flash_io0_oeb 30.62fF
C3565 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<15> 0.05fF
C3566 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<10> 11.12fF
C3567 LOGIC1_3V_2|Q LOGIC1_3V_1|Q 0.58fF
C3568 BU_3VX2_9|A LS_3VX2_3|Q 1.82fF
C3569 BU_3VX2_16|A BU_3VX2_28|A 1.73fF
C3570 BU_3VX2_29|A BU_3VX2_28|A 90.58fF
C3571 AMUX4_3V_0|AIN1 BU_3VX2_47|A 0.02fF
C3572 LS_3VX2_12|A BU_3VX2_60|Q 0.01fF
C3573 LOGIC0_3V_4|Q raven_soc_0|flash_clk 0.22fF
C3574 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<9> 0.75fF
C3575 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pullup<14> 0.01fF
C3576 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<5> 1.02fF
C3577 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<14> 0.03fF
C3578 LS_3VX2_13|A BU_3VX2_59|Q 0.01fF
C3579 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_11|PO 0.04fF
C3580 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<6> 0.01fF
C3581 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<29> 37.35fF
C3582 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<5> 0.01fF
C3583 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<7> 0.01fF
C3584 BU_3VX2_1|Q AMUX4_3V_4|SEL[1] 1.69fF
C3585 BU_3VX2_66|Q BU_3VX2_22|Q 2.26fF
C3586 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<19> 7.18fF
C3587 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<31> 3.41fF
C3588 BU_3VX2_38|Q BU_3VX2_2|Q 21.82fF
C3589 BU_3VX2_12|Q BU_3VX2_8|Q 13.05fF
C3590 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<25> 0.63fF
C3591 BU_3VX2_2|Q BU_3VX2_67|Q 1.34fF
C3592 BU_3VX2_15|Q BU_3VX2_17|Q 24.30fF
C3593 BU_3VX2_12|Q BU_3VX2_21|Q 5.75fF
C3594 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<17> 1.00fF
C3595 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<21> 10.23fF
C3596 LS_3VX2_2|A AMUX4_3V_3|SEL[0] 1.54fF
C3597 BU_3VX2_38|Q BU_3VX2_10|Q 2.81fF
C3598 BU_3VX2_67|Q BU_3VX2_10|Q 0.58fF
C3599 raven_soc_0|gpio_in<8> vdd 1.78fF
C3600 BU_3VX2_9|Q BU_3VX2_17|Q 4.16fF
C3601 BU_3VX2_22|Q BU_3VX2_20|Q 21.30fF
C3602 raven_soc_0|ext_clk BU_3VX2_23|Q 0.01fF
C3603 BU_3VX2_60|A vdd 0.07fF
C3604 VDD3V3 BU_3VX2_28|Q 2.22fF
C3605 BU_3VX2_24|A BU_3VX2_14|A 2.02fF
C3606 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<4> 0.01fF
C3607 raven_padframe_0|BBC4F_1|VDDO raven_padframe_0|BBC4F_1|GNDO 2.28fF
C3608 BU_3VX2_21|A BU_3VX2_13|A 2.03fF
C3609 BU_3VX2_37|A BU_3VX2_28|A 0.01fF
C3610 LS_3VX2_10|Q LS_3VX2_14|Q 0.74fF
C3611 raven_padframe_0|aregc01_3v3_1|m4_0_29333# raven_padframe_0|aregc01_3v3_1|m4_0_28769# 0.03fF
C3612 raven_padframe_0|APR00DF_2|VDDR raven_padframe_0|APR00DF_2|GNDO 0.13fF
C3613 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<5> 2.45fF
C3614 raven_padframe_0|axtoc02_3v3_0|m4_0_30133# raven_padframe_0|axtoc02_3v3_0|m4_0_29333# 0.17fF
C3615 raven_soc_0|gpio_out<3> BU_3VX2_0|Q 0.01fF
C3616 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<9> 17.02fF
C3617 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<8> 0.01fF
C3618 BU_3VX2_63|Q raven_soc_0|gpio_pullup<11> 0.01fF
C3619 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<10> 22.91fF
C3620 BU_3VX2_10|A VDD3V3 0.21fF
C3621 raven_soc_0|gpio_out<4> raven_soc_0|ext_clk 0.01fF
C3622 LS_3VX2_4|A VDD3V3 0.53fF
C3623 LS_3VX2_7|A BU_3VX2_48|Q 0.03fF
C3624 raven_soc_0|gpio_pulldown<12> VDD3V3 0.07fF
C3625 BU_3VX2_1|Q raven_soc_0|flash_io2_oeb 0.01fF
C3626 raven_soc_0|gpio_pulldown<3> apllc03_1v8_0|CLK 0.01fF
C3627 raven_soc_0|gpio_pullup<13> vdd 0.22fF
C3628 BU_3VX2_73|Q BU_3VX2_47|Q 8.66fF
C3629 LOGIC0_3V_0|Q LOGIC0_3V_3|Q 6.00fF
C3630 raven_spi_0|CSB raven_soc_0|gpio_pulldown<15> 1.51fF
C3631 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_out<3> 1.68fF
C3632 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<13> 1.86fF
C3633 BU_3VX2_0|A VDD3V3 0.86fF
C3634 IN_3VX2_1|Q BU_3VX2_50|Q 0.49fF
C3635 VDD raven_padframe_0|FILLER20F_7|VDDR 0.71fF
C3636 LS_3VX2_7|A raven_soc_0|ser_tx 0.01fF
C3637 LS_3VX2_24|A AMUX4_3V_1|SEL[1] 0.02fF
C3638 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<8> 0.50fF
C3639 AMUX4_3V_4|AIN1 comp_inp 57.35fF
C3640 BU_3VX2_0|Q raven_soc_0|ram_wdata<26> 0.02fF
C3641 BU_3VX2_26|A vdd 0.06fF
C3642 VDD raven_padframe_0|axtoc02_3v3_0|m4_0_31172# 0.25fF
C3643 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<15> 0.72fF
C3644 raven_soc_0|flash_io1_oeb raven_soc_0|flash_clk 136.26fF
C3645 raven_padframe_0|BBC4F_0|VDDO raven_padframe_0|BBC4F_0|GNDO 2.28fF
C3646 raven_padframe_0|BBCUD4F_4|GNDR raven_padframe_0|BBCUD4F_4|GNDO 0.81fF
C3647 raven_soc_0|gpio_in<1> apllc03_1v8_0|CLK 0.02fF
C3648 LS_3VX2_7|A LS_3VX2_24|A 12.48fF
C3649 BU_3VX2_23|A raven_soc_0|flash_io2_do 0.01fF
C3650 BU_3VX2_9|A raven_soc_0|flash_io1_oeb 0.01fF
C3651 BU_3VX2_19|A raven_soc_0|flash_io0_do 0.01fF
C3652 raven_padframe_0|ICFC_1|VDD3 raven_padframe_0|ICFC_1|GNDO 0.07fF
C3653 BU_3VX2_31|A raven_soc_0|gpio_out<10> 0.01fF
C3654 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<13> 0.01fF
C3655 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<8> 0.35fF
C3656 AMUX4_3V_4|AIN1 AMUX4_3V_4|SEL[0] 0.02fF
C3657 IN_3VX2_1|A BU_3VX2_29|Q 101.96fF
C3658 BU_3VX2_11|A vdd 0.06fF
C3659 raven_padframe_0|BBCUD4F_12|VDDR raven_padframe_0|BBCUD4F_12|GNDO 0.13fF
C3660 raven_soc_0|ser_rx BU_3VX2_59|Q 2.51fF
C3661 raven_soc_0|gpio_outenb<5> apllc03_1v8_0|CLK 0.01fF
C3662 raven_soc_0|gpio_out<5> vdd 0.18fF
C3663 raven_soc_0|gpio_outenb<11> BU_3VX2_24|Q 0.01fF
C3664 raven_soc_0|gpio_outenb<14> BU_3VX2_26|Q 0.01fF
C3665 raven_soc_0|gpio_pullup<12> BU_3VX2_27|Q 0.01fF
C3666 raven_soc_0|gpio_outenb<10> BU_3VX2_23|Q 0.01fF
C3667 raven_soc_0|gpio_outenb<12> BU_3VX2_25|Q 0.01fF
C3668 LS_3VX2_3|Q BU_3VX2_28|A 0.01fF
C3669 BU_3VX2_1|A BU_3VX2_64|A 0.59fF
C3670 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<10> 0.09fF
C3671 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<3> 0.72fF
C3672 BU_3VX2_25|A raven_soc_0|flash_io0_oeb 3.66fF
C3673 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<6> 0.01fF
C3674 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<8> 6.42fF
C3675 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<4> 0.01fF
C3676 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<14> 0.15fF
C3677 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<10> 5.84fF
C3678 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<10> 1.80fF
C3679 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<15> 16.81fF
C3680 raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<11> 2.56fF
C3681 BU_3VX2_40|Q raven_soc_0|flash_io3_do 0.01fF
C3682 VDD3V3 comp_inp 8.41fF
C3683 BU_3VX2_61|A LS_3VX2_17|Q 0.82fF
C3684 BU_3VX2_60|A BU_3VX2_62|A 0.73fF
C3685 LS_3VX2_15|Q LS_3VX2_16|Q 16.46fF
C3686 VDD3V3 BU_3VX2_44|Q 1.43fF
C3687 LS_3VX2_9|A LS_3VX2_6|A 33.02fF
C3688 BU_3VX2_16|A BU_3VX2_14|A 13.56fF
C3689 BU_3VX2_40|A BU_3VX2_11|A 1.01fF
C3690 raven_padframe_0|FILLER20F_4|GNDR raven_padframe_0|FILLER20F_4|VDDO 0.09fF
C3691 BU_3VX2_18|A raven_soc_0|flash_csb 0.01fF
C3692 BU_3VX2_29|A BU_3VX2_14|A 0.01fF
C3693 raven_padframe_0|aregc01_3v3_0|m4_0_29057# raven_padframe_0|aregc01_3v3_0|m4_0_28769# 0.11fF
C3694 raven_padframe_0|APR00DF_0|GNDR raven_padframe_0|APR00DF_0|VDDO 0.09fF
C3695 BU_3VX2_31|A raven_soc_0|gpio_out<9> 0.01fF
C3696 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<5> 0.02fF
C3697 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<4> 0.84fF
C3698 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<9> 0.34fF
C3699 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<11> 0.19fF
C3700 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<6> 1.95fF
C3701 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<28> 0.68fF
C3702 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<20> 0.08fF
C3703 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<23> 0.05fF
C3704 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<11> 0.01fF
C3705 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<11> 7.13fF
C3706 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<8> 11.64fF
C3707 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<12> 8.33fF
C3708 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_out<15> 0.02fF
C3709 raven_soc_0|gpio_out<14> BU_3VX2_40|Q 0.01fF
C3710 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<10> 0.02fF
C3711 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<2> 0.14fF
C3712 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<1> 0.23fF
C3713 raven_soc_0|ram_wdata<10> vdd 0.67fF
C3714 AMUX4_3V_4|SEL[0] VDD3V3 0.73fF
C3715 LS_3VX2_21|A BU_3VX2_49|Q 20.27fF
C3716 LS_3VX2_27|A BU_3VX2_51|Q 28.56fF
C3717 AMUX4_3V_0|SEL[1] LS_3VX2_27|A 0.52fF
C3718 raven_soc_0|gpio_in<8> raven_padframe_0|BBCUD4F_8|PO 0.04fF
C3719 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<4> 1.97fF
C3720 raven_padframe_0|VDDPADF_0|VDDR raven_padframe_0|VDDPADF_0|VDDO 0.06fF
C3721 BU_3VX2_37|A BU_3VX2_14|A 0.94fF
C3722 LS_3VX2_11|Q LS_3VX2_24|Q 0.01fF
C3723 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<0> 128.76fF
C3724 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<12> 0.35fF
C3725 LS_3VX2_13|A AMUX2_3V_0|SEL 53.02fF
C3726 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<8> 0.01fF
C3727 LS_3VX2_14|A BU_3VX2_54|Q 0.02fF
C3728 AMUX4_3V_4|AIN1 vdd 4.84fF
C3729 BU_3VX2_0|Q BU_3VX2_22|Q 0.01fF
C3730 VDD raven_padframe_0|CORNERESDF_1|GNDR 0.16fF
C3731 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_outenb<9> 1.56fF
C3732 raven_soc_0|gpio_out<10> raven_soc_0|gpio_out<8> 7.64fF
C3733 raven_soc_0|gpio_pulldown<7> BU_3VX2_71|Q 0.38fF
C3734 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<5> 0.09fF
C3735 raven_soc_0|ram_rdata<14> raven_soc_0|ram_addr<4> 1.38fF
C3736 raven_soc_0|ram_rdata<24> raven_soc_0|ram_addr<3> 7.05fF
C3737 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<6> 0.08fF
C3738 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<7> 0.30fF
C3739 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<8> 0.12fF
C3740 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<9> 7.63fF
C3741 raven_soc_0|ram_rdata<21> raven_soc_0|ram_addr<2> 4.07fF
C3742 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<30> 0.45fF
C3743 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<20> 0.01fF
C3744 BU_3VX2_24|A raven_soc_0|flash_io1_do 0.01fF
C3745 LOGIC0_3V_0|Q VDD3V3 0.28fF
C3746 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<7> 2.62fF
C3747 BU_3VX2_3|A raven_soc_0|flash_io3_do 0.01fF
C3748 BU_3VX2_15|A raven_soc_0|flash_io3_do 0.01fF
C3749 IN_3VX2_1|A raven_soc_0|flash_io2_do 4.64fF
C3750 BU_3VX2_67|A BU_3VX2_65|Q 0.03fF
C3751 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<14> 0.03fF
C3752 BU_3VX2_28|A raven_soc_0|flash_io1_oeb 6.83fF
C3753 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<11> 2.59fF
C3754 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<9> 7.59fF
C3755 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<13> 68.63fF
C3756 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<10> 0.44fF
C3757 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<6> 6.35fF
C3758 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<7> 0.02fF
C3759 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<15> 0.02fF
C3760 raven_padframe_0|ICFC_1|VDD3 raven_padframe_0|ICFC_1|VDDR 0.71fF
C3761 BU_3VX2_20|A BU_3VX2_18|A 12.50fF
C3762 LS_3VX2_13|Q LS_3VX2_5|Q 0.75fF
C3763 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<8> 0.01fF
C3764 raven_spi_0|SDO raven_soc_0|gpio_pullup<15> 1.13fF
C3765 BU_3VX2_1|A BU_3VX2_66|A 0.52fF
C3766 LS_3VX2_12|A BU_3VX2_62|Q 0.01fF
C3767 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<6> 0.01fF
C3768 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<8> 0.01fF
C3769 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_outenb<13> 31.50fF
C3770 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<10> 0.78fF
C3771 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<8> 0.98fF
C3772 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<8> 11.03fF
C3773 raven_soc_0|gpio_out<5> raven_soc_0|gpio_outenb<9> 0.01fF
C3774 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<5> 0.01fF
C3775 raven_soc_0|ram_wenb raven_soc_0|ram_addr<0> 0.01fF
C3776 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<14> 0.02fF
C3777 LS_3VX2_13|A BU_3VX2_61|Q 0.01fF
C3778 BU_3VX2_19|Q BU_3VX2_12|Q 6.23fF
C3779 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<25> 160.41fF
C3780 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<2> 0.47fF
C3781 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<29> 0.11fF
C3782 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<15> 0.01fF
C3783 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<17> 133.81fF
C3784 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<21> 3.32fF
C3785 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<14> 102.16fF
C3786 BU_3VX2_13|Q BU_3VX2_69|Q 22.88fF
C3787 BU_3VX2_21|Q BU_3VX2_5|Q 0.15fF
C3788 BU_3VX2_12|Q BU_3VX2_18|Q 78.41fF
C3789 BU_3VX2_66|Q BU_3VX2_31|Q 0.45fF
C3790 BU_3VX2_6|Q BU_3VX2_7|Q 69.85fF
C3791 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<19> 1.41fF
C3792 BU_3VX2_16|Q BU_3VX2_22|Q 5.66fF
C3793 raven_soc_0|ram_wdata<8> raven_soc_0|ram_rdata<2> 0.01fF
C3794 BU_3VX2_30|Q BU_3VX2_22|Q 6.22fF
C3795 BU_3VX2_31|Q BU_3VX2_20|Q 22.68fF
C3796 BU_3VX2_5|Q BU_3VX2_8|Q 18.03fF
C3797 BU_3VX2_65|Q BU_3VX2_10|Q 0.93fF
C3798 BU_3VX2_33|Q BU_3VX2_67|Q 0.54fF
C3799 VDD3V3 vdd 193.03fF
C3800 BU_3VX2_56|Q BU_3VX2_54|Q 80.37fF
C3801 LS_3VX2_7|Q LS_3VX2_10|Q 2.22fF
C3802 LS_3VX2_11|Q LS_3VX2_6|Q 12.33fF
C3803 LS_3VX2_12|A LS_3VX2_5|A 20.45fF
C3804 LOGIC1_3V_3|Q LOGIC0_3V_2|Q 0.21fF
C3805 raven_padframe_0|BBCUD4F_10|GNDR raven_padframe_0|BBCUD4F_10|VDDO 0.09fF
C3806 BU_3VX2_37|A LS_3VX2_3|A 0.49fF
C3807 LS_3VX2_3|Q BU_3VX2_14|A 0.01fF
C3808 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<7> 0.01fF
C3809 BU_3VX2_69|A BU_3VX2_36|A 1.93fF
C3810 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<4> 0.01fF
C3811 AMUX2_3V_0|SEL raven_soc_0|ser_rx 0.01fF
C3812 raven_soc_0|flash_io1_oeb BU_3VX2_33|Q 0.01fF
C3813 LS_3VX2_8|Q LS_3VX2_11|Q 2.80fF
C3814 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<7> 0.66fF
C3815 BU_3VX2_71|A raven_soc_0|flash_csb 0.01fF
C3816 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<15> 0.01fF
C3817 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<6> 1.34fF
C3818 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<12> 0.65fF
C3819 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<6> 0.36fF
C3820 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<8> 0.01fF
C3821 IN_3VX2_1|Q BU_3VX2_48|Q 0.61fF
C3822 BU_3VX2_40|A VDD3V3 1.17fF
C3823 VDD raven_padframe_0|CORNERESDF_2|GNDR 0.16fF
C3824 raven_padframe_0|FILLER20F_8|VDDR raven_padframe_0|FILLER20F_8|VDDO 0.06fF
C3825 VDD raven_padframe_0|FILLER40F_0|GNDR 0.16fF
C3826 raven_soc_0|gpio_pulldown<1> BU_3VX2_40|Q 0.03fF
C3827 BU_3VX2_31|A raven_soc_0|ext_clk 0.16fF
C3828 BU_3VX2_0|Q raven_soc_0|ram_wdata<28> 0.02fF
C3829 raven_soc_0|gpio_in<2> VDD3V3 3.00fF
C3830 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<17> 0.09fF
C3831 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<31> 14.03fF
C3832 raven_soc_0|ram_addr<4> raven_soc_0|ram_addr<0> 16.59fF
C3833 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<27> 0.12fF
C3834 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<15> 0.07fF
C3835 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<13> 10.39fF
C3836 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<1> 0.01fF
C3837 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<16> 0.01fF
C3838 BU_3VX2_59|Q BU_3VX2_72|Q 0.17fF
C3839 raven_soc_0|gpio_out<1> IN_3VX2_1|A 0.01fF
C3840 BU_3VX2_19|A raven_soc_0|flash_io1_di 0.01fF
C3841 BU_3VX2_16|A raven_soc_0|flash_io1_do 0.06fF
C3842 BU_3VX2_4|A raven_soc_0|flash_io0_oeb 0.01fF
C3843 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<7> 0.01fF
C3844 raven_padframe_0|ICF_2|VDDR raven_padframe_0|ICF_2|GNDR 0.68fF
C3845 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<5> 1.63fF
C3846 BU_3VX2_29|A raven_soc_0|flash_io1_do 4.61fF
C3847 BU_3VX2_64|A BU_3VX2_1|Q 0.03fF
C3848 raven_soc_0|gpio_pullup<10> BU_3VX2_23|Q 0.01fF
C3849 raven_soc_0|gpio_outenb<6> vdd 0.34fF
C3850 raven_soc_0|gpio_pullup<15> BU_3VX2_26|Q 0.01fF
C3851 raven_soc_0|gpio_pullup<11> BU_3VX2_24|Q 0.01fF
C3852 raven_soc_0|gpio_pullup<8> BU_3VX2_28|Q 0.01fF
C3853 raven_soc_0|gpio_outenb<0> BU_3VX2_27|Q 0.04fF
C3854 raven_soc_0|gpio_pullup<12> BU_3VX2_25|Q 0.01fF
C3855 raven_soc_0|ser_rx BU_3VX2_61|Q 3.31fF
C3856 raven_soc_0|gpio_pullup<7> apllc03_1v8_0|CLK 0.01fF
C3857 LS_3VX2_3|Q LS_3VX2_3|A 0.03fF
C3858 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<13> 0.01fF
C3859 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<10> 0.01fF
C3860 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<8> 0.01fF
C3861 BU_3VX2_35|A raven_soc_0|flash_io3_oeb 0.01fF
C3862 BU_3VX2_37|A raven_soc_0|flash_io1_do 0.01fF
C3863 AMUX4_3V_4|AOUT raven_soc_0|flash_io0_oeb 3.59fF
C3864 BU_3VX2_25|A raven_soc_0|flash_io2_do 0.01fF
C3865 BU_3VX2_14|A raven_soc_0|flash_io1_oeb 0.01fF
C3866 LOGIC0_3V_4|Q raven_padframe_0|ICFC_0|PO 0.04fF
C3867 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<13> 30.15fF
C3868 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<12> 3.02fF
C3869 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<7> 0.69fF
C3870 raven_soc_0|gpio_in<11> VDD3V3 0.07fF
C3871 BU_3VX2_53|A LS_3VX2_15|Q 0.15fF
C3872 BU_3VX2_52|A LS_3VX2_16|Q 0.11fF
C3873 BU_3VX2_57|A BU_3VX2_58|A 7.98fF
C3874 BU_3VX2_56|A BU_3VX2_59|A 1.28fF
C3875 BU_3VX2_55|A BU_3VX2_60|A 0.59fF
C3876 BU_3VX2_54|A BU_3VX2_61|A 0.32fF
C3877 VDD3V3 BU_3VX2_62|A 0.08fF
C3878 LS_3VX2_20|A BU_3VX2_43|Q 8.91fF
C3879 BU_3VX2_3|A BU_3VX2_8|A 2.37fF
C3880 BU_3VX2_2|A BU_3VX2_35|A 6.02fF
C3881 BU_3VX2_8|A BU_3VX2_15|A 1.72fF
C3882 BU_3VX2_20|A BU_3VX2_71|A 0.01fF
C3883 LS_3VX2_19|Q aopac01_3v3_0|IB 0.66fF
C3884 raven_spi_0|SDI BU_3VX2_33|A 70.96fF
C3885 BU_3VX2_31|A raven_soc_0|gpio_outenb<10> 0.01fF
C3886 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<6> 0.01fF
C3887 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<2> 4.18fF
C3888 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<9> 0.01fF
C3889 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<6> 25.24fF
C3890 raven_soc_0|gpio_out<8> raven_soc_0|ext_clk 0.01fF
C3891 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<13> 0.02fF
C3892 raven_soc_0|gpio_outenb<9> VDD3V3 0.07fF
C3893 BU_3VX2_21|Q BU_3VX2_28|Q 6.09fF
C3894 BU_3VX2_12|Q BU_3VX2_27|Q 4.67fF
C3895 BU_3VX2_8|Q BU_3VX2_28|Q 5.55fF
C3896 BU_3VX2_13|Q BU_3VX2_29|Q 0.09fF
C3897 BU_3VX2_66|Q apllc03_1v8_0|CLK 0.94fF
C3898 BU_3VX2_20|Q apllc03_1v8_0|CLK 0.01fF
C3899 LS_3VX2_27|A BU_3VX2_49|Q 15.76fF
C3900 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<15> 0.01fF
C3901 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<12> 0.01fF
C3902 BU_3VX2_10|A BU_3VX2_8|Q 0.03fF
C3903 LS_3VX2_14|A BU_3VX2_56|Q 0.05fF
C3904 BU_3VX2_0|Q BU_3VX2_31|Q 0.25fF
C3905 adc_high AMUX4_3V_4|AIN2 2.02fF
C3906 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<23> 0.02fF
C3907 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<4> 9.60fF
C3908 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<18> 27.86fF
C3909 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<24> 0.44fF
C3910 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<14> 2.78fF
C3911 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_out<10> 0.02fF
C3912 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pullup<14> 0.02fF
C3913 AMUX4_3V_1|SEL[0] BU_3VX2_59|Q 12.79fF
C3914 raven_soc_0|flash_io0_do BU_3VX2_27|Q 0.01fF
C3915 raven_soc_0|ram_rdata<28> apllc03_1v8_0|CLK 0.01fF
C3916 raven_padframe_0|axtoc02_3v3_0|m4_55000_28769# raven_padframe_0|axtoc02_3v3_0|GNDO 0.07fF
C3917 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<15> 1.49fF
C3918 raven_soc_0|gpio_out<0> BU_3VX2_40|Q 0.02fF
C3919 BU_3VX2_22|A raven_soc_0|ext_clk 0.01fF
C3920 LS_3VX2_3|Q raven_soc_0|flash_io1_do 0.01fF
C3921 raven_padframe_0|ICF_1|VDDR raven_padframe_0|ICF_1|GNDO 0.13fF
C3922 raven_soc_0|gpio_out<6> raven_soc_0|ext_clk 0.01fF
C3923 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<13> 12.83fF
C3924 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<6> 0.01fF
C3925 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<8> 0.39fF
C3926 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<7> 0.34fF
C3927 LS_3VX2_3|A raven_soc_0|flash_io1_oeb 0.62fF
C3928 raven_soc_0|gpio_out<12> BU_3VX2_40|Q 0.01fF
C3929 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pullup<5> 1.53fF
C3930 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<11> 0.02fF
C3931 BU_3VX2_0|Q raven_soc_0|flash_io3_oeb 0.01fF
C3932 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<15> 0.02fF
C3933 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<19> 6.07fF
C3934 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<0> 1.26fF
C3935 BU_3VX2_10|A BU_3VX2_19|A 1.41fF
C3936 LOGIC0_3V_4|Q raven_soc_0|flash_io1_do 0.01fF
C3937 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<9> 1.40fF
C3938 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<8> 3.81fF
C3939 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<13> 9.06fF
C3940 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<10> 12.26fF
C3941 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pullup<13> 75.88fF
C3942 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<14> 0.02fF
C3943 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<5> 0.01fF
C3944 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<8> 24.63fF
C3945 raven_soc_0|ram_wenb raven_soc_0|ram_addr<9> 0.01fF
C3946 raven_soc_0|gpio_pullup<4> BU_3VX2_71|Q 0.01fF
C3947 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pulldown<6> 1.83fF
C3948 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<6> 0.01fF
C3949 raven_soc_0|gpio_pulldown<15> apllc03_1v8_0|CLK 1.20fF
C3950 LS_3VX2_13|A LS_3VX2_15|A 0.02fF
C3951 raven_soc_0|gpio_pulldown<14> BU_3VX2_27|Q 0.01fF
C3952 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<18> 48.60fF
C3953 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<3> 0.10fF
C3954 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<26> 0.25fF
C3955 raven_spi_0|CSB raven_spi_0|SDO 100.76fF
C3956 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<1> 0.01fF
C3957 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<25> 0.01fF
C3958 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<15> 13.71fF
C3959 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<12> 0.02fF
C3960 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<14> 9.49fF
C3961 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<8> 4.99fF
C3962 BU_3VX2_35|Q BU_3VX2_6|Q 3.83fF
C3963 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<13> 3.90fF
C3964 raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<8> 10.28fF
C3965 BU_3VX2_19|Q BU_3VX2_5|Q 0.22fF
C3966 BU_3VX2_31|Q BU_3VX2_30|Q 58.57fF
C3967 BU_3VX2_68|Q BU_3VX2_9|Q 0.99fF
C3968 BU_3VX2_5|Q BU_3VX2_18|Q 2.39fF
C3969 raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<14> 1.50fF
C3970 BU_3VX2_35|Q BU_3VX2_7|Q 3.25fF
C3971 BU_3VX2_65|Q BU_3VX2_33|Q 0.52fF
C3972 raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<13> 1.39fF
C3973 BU_3VX2_57|Q BU_3VX2_55|Q 82.02fF
C3974 LS_3VX2_20|A BU_3VX2_50|Q 56.25fF
C3975 BU_3VX2_19|A BU_3VX2_0|A 0.01fF
C3976 LS_3VX2_10|Q LS_3VX2_4|Q 1.33fF
C3977 BU_3VX2_73|A LS_3VX2_24|Q 1.79fF
C3978 raven_soc_0|gpio_outenb<4> BU_3VX2_0|Q 0.26fF
C3979 raven_soc_0|ram_wdata<25> vdd 1.09fF
C3980 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<13> 0.15fF
C3981 BU_3VX2_24|A raven_soc_0|flash_csb 4.56fF
C3982 vdd raven_padframe_0|VDDPADF_1|GNDR 0.16fF
C3983 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<7> 0.01fF
C3984 LS_3VX2_9|Q LS_3VX2_6|A 0.18fF
C3985 IN_3VX2_1|A raven_soc_0|gpio_out<11> 0.01fF
C3986 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<13> 0.23fF
C3987 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<5> 0.13fF
C3988 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<9> 5.08fF
C3989 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<6> 0.01fF
C3990 raven_soc_0|gpio_outenb<2> BU_3VX2_63|Q 0.01fF
C3991 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<11> 0.01fF
C3992 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<12> 0.02fF
C3993 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<7> 0.01fF
C3994 raven_soc_0|gpio_pulldown<2> raven_soc_0|ext_clk 0.01fF
C3995 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io3_di 46.90fF
C3996 BU_3VX2_2|Q BU_3VX2_36|Q 2.18fF
C3997 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<31> 3.81fF
C3998 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io0_do 139.76fF
C3999 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<17> 124.24fF
C4000 raven_soc_0|ram_addr<9> raven_soc_0|ram_addr<4> 7.95fF
C4001 raven_soc_0|flash_io1_do raven_soc_0|flash_io1_oeb 61.93fF
C4002 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<19> 17.58fF
C4003 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<13> 83.06fF
C4004 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<10> 0.53fF
C4005 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<26> 0.37fF
C4006 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<1> 7.10fF
C4007 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<15> 4.36fF
C4008 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<25> 2.30fF
C4009 raven_soc_0|ram_rdata<5> raven_soc_0|ram_addr<0> 0.09fF
C4010 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<24> 0.01fF
C4011 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<29> 0.01fF
C4012 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<27> 0.01fF
C4013 raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<2> 8.45fF
C4014 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<22> 0.01fF
C4015 BU_3VX2_36|Q BU_3VX2_10|Q 1.06fF
C4016 LS_3VX2_17|A BU_3VX2_59|Q 17.33fF
C4017 BU_3VX2_45|A BU_3VX2_43|Q 0.03fF
C4018 BU_3VX2_43|Q BU_3VX2_47|Q 25.76fF
C4019 BU_3VX2_44|Q adc0_data<5> 47.55fF
C4020 BU_3VX2_45|Q BU_3VX2_46|Q 216.68fF
C4021 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<3> 0.01fF
C4022 BU_3VX2_6|A raven_soc_0|flash_io0_do 0.02fF
C4023 BU_3VX2_21|A raven_soc_0|ext_clk 0.17fF
C4024 BU_3VX2_2|A raven_soc_0|flash_io3_di 0.02fF
C4025 BU_3VX2_4|A raven_soc_0|flash_io2_do 0.01fF
C4026 raven_soc_0|gpio_pullup<2> VDD3V3 4.87fF
C4027 BU_3VX2_38|A raven_soc_0|flash_io2_di 0.01fF
C4028 LS_3VX2_5|Q LS_3VX2_19|A 0.01fF
C4029 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<6> 0.60fF
C4030 IN_3VX2_1|A AMUX4_3V_4|AIN2 3.77fF
C4031 raven_padframe_0|BBCUD4F_13|VDDR raven_padframe_0|BBCUD4F_13|GNDO 0.13fF
C4032 raven_soc_0|gpio_pullup<8> vdd 0.23fF
C4033 BU_3VX2_0|Q apllc03_1v8_0|CLK 110.70fF
C4034 VDD raven_padframe_0|BBCUD4F_2|GNDR 0.16fF
C4035 raven_soc_0|ser_rx LS_3VX2_15|A 4.24fF
C4036 raven_soc_0|gpio_pulldown<10> BU_3VX2_27|Q 0.01fF
C4037 raven_soc_0|gpio_outenb<0> BU_3VX2_25|Q 0.01fF
C4038 BU_3VX2_71|Q raven_soc_0|flash_clk 0.33fF
C4039 raven_soc_0|gpio_in<3> raven_padframe_0|BBCUD4F_3|PO 0.04fF
C4040 LS_3VX2_13|Q LS_3VX2_12|Q 5.59fF
C4041 BU_3VX2_7|A BU_3VX2_26|A 0.01fF
C4042 raven_soc_0|gpio_pulldown<13> LS_3VX2_3|A 0.01fF
C4043 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<4> 1.19fF
C4044 BU_3VX2_70|A BU_3VX2_0|Q 1.34fF
C4045 VDD raven_padframe_0|BBCUD4F_6|GNDR 0.16fF
C4046 AMUX2_3V_0|SEL AMUX4_3V_1|SEL[0] 8.61fF
C4047 raven_soc_0|gpio_pulldown<0> apllc03_1v8_0|CLK 0.22fF
C4048 LS_3VX2_13|A AMUX4_3V_1|SEL[1] 8.17fF
C4049 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<15> 0.02fF
C4050 BU_3VX2_24|A BU_3VX2_20|A 5.65fF
C4051 BU_3VX2_40|Q raven_soc_0|gpio_pullup<5> 0.01fF
C4052 BU_3VX2_52|A BU_3VX2_53|A 13.29fF
C4053 VDD3V3 BU_3VX2_55|A 0.05fF
C4054 raven_padframe_0|POWERCUTVDD3FC_0|VDDO raven_padframe_0|POWERCUTVDD3FC_0|GNDO 2.22fF
C4055 BU_3VX2_7|A BU_3VX2_11|A 3.06fF
C4056 LS_3VX2_5|Q adc_low 0.12fF
C4057 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<9> 0.06fF
C4058 LS_3VX2_7|A LS_3VX2_13|A 32.13fF
C4059 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<4> 4.98fF
C4060 LS_3VX2_24|Q LS_3VX2_4|A 0.16fF
C4061 BU_3VX2_31|A raven_soc_0|gpio_pullup<10> 0.01fF
C4062 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<8> 0.01fF
C4063 raven_soc_0|gpio_pullup<1> LS_3VX2_3|A 0.13fF
C4064 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<13> 0.30fF
C4065 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<8> 0.01fF
C4066 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<5> 0.01fF
C4067 raven_soc_0|flash_io3_oeb raven_soc_0|irq_pin 0.01fF
C4068 raven_soc_0|gpio_pulldown<6> raven_soc_0|ext_clk 0.01fF
C4069 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<9> 3.74fF
C4070 BU_3VX2_5|Q BU_3VX2_27|Q 2.23fF
C4071 BU_3VX2_9|Q BU_3VX2_24|Q 1.54fF
C4072 BU_3VX2_12|Q BU_3VX2_25|Q 17.68fF
C4073 BU_3VX2_18|Q BU_3VX2_28|Q 6.25fF
C4074 BU_3VX2_8|Q vdd 1.15fF
C4075 BU_3VX2_21|Q vdd 0.98fF
C4076 BU_3VX2_19|Q BU_3VX2_28|Q 17.88fF
C4077 BU_3VX2_22|Q BU_3VX2_26|Q 9.80fF
C4078 BU_3VX2_7|Q BU_3VX2_23|Q 2.86fF
C4079 BU_3VX2_69|Q BU_3VX2_29|Q 0.48fF
C4080 LS_3VX2_16|A BU_3VX2_55|Q 11.14fF
C4081 AMUX4_3V_0|SEL[1] BU_3VX2_53|Q 0.14fF
C4082 BU_3VX2_6|Q BU_3VX2_23|Q 0.59fF
C4083 BU_3VX2_33|Q BU_3VX2_72|Q 0.14fF
C4084 BU_3VX2_15|Q BU_3VX2_24|Q 3.96fF
C4085 BU_3VX2_16|Q apllc03_1v8_0|CLK 0.01fF
C4086 BU_3VX2_30|Q apllc03_1v8_0|CLK 3.34fF
C4087 LS_3VX2_12|A LS_3VX2_11|A 74.97fF
C4088 raven_padframe_0|ICFC_2|VDD3 LOGIC0_3V_4|Q 0.04fF
C4089 LS_3VX2_8|Q LS_3VX2_8|A 0.05fF
C4090 LS_3VX2_11|Q LS_3VX2_14|Q 0.47fF
C4091 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<6> 2.03fF
C4092 BU_3VX2_16|A raven_soc_0|flash_csb 0.01fF
C4093 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<2> 113.68fF
C4094 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<12> 0.01fF
C4095 BU_3VX2_29|A raven_soc_0|flash_csb 17.91fF
C4096 AMUX4_3V_3|SEL[1] BU_3VX2_14|Q 1.29fF
C4097 raven_soc_0|ram_rdata<1> raven_soc_0|ram_rdata<15> 0.04fF
C4098 raven_soc_0|ram_rdata<13> raven_soc_0|ram_addr<0> 0.01fF
C4099 raven_soc_0|ram_wdata<31> raven_soc_0|ram_rdata<16> 0.01fF
C4100 AMUX4_3V_1|SEL[0] BU_3VX2_61|Q 9.62fF
C4101 raven_soc_0|flash_io0_oeb BU_3VX2_29|Q 11.03fF
C4102 raven_soc_0|flash_io3_di apllc03_1v8_0|CLK 17.46fF
C4103 raven_soc_0|flash_io1_di BU_3VX2_27|Q 0.01fF
C4104 LS_3VX2_15|Q BU_3VX2_58|Q 0.11fF
C4105 raven_soc_0|flash_io0_do BU_3VX2_25|Q 0.01fF
C4106 raven_soc_0|flash_io2_di BU_3VX2_23|Q 0.01fF
C4107 BU_3VX2_47|Q BU_3VX2_50|Q 45.57fF
C4108 adc0_data<5> vdd 1.83fF
C4109 BU_3VX2_37|A raven_soc_0|flash_csb 0.01fF
C4110 markings_0|manufacturer_0|_alphabet_S_1|m2_32_224# markings_0|manufacturer_0|_alphabet_S_0|m2_32_224# 0.45fF
C4111 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<14> 0.26fF
C4112 BU_3VX2_63|A raven_soc_0|flash_io3_oeb 0.01fF
C4113 BU_3VX2_19|A vdd 0.06fF
C4114 LS_3VX2_6|A BU_3VX2_73|Q 8.66fF
C4115 IN_3VX2_1|A raven_soc_0|gpio_in<12> 0.01fF
C4116 raven_soc_0|gpio_outenb<12> BU_3VX2_40|Q 0.01fF
C4117 BU_3VX2_69|A VDD3V3 0.02fF
C4118 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<8> 0.01fF
C4119 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<7> 0.01fF
C4120 raven_soc_0|gpio_outenb<14> VDD3V3 0.07fF
C4121 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<6> 0.01fF
C4122 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pullup<5> 1.78fF
C4123 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<11> 3.70fF
C4124 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<15> 0.02fF
C4125 raven_soc_0|gpio_outenb<11> raven_soc_0|ext_clk 0.01fF
C4126 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<23> 0.65fF
C4127 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<20> 0.63fF
C4128 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<11> 23.72fF
C4129 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<19> 6.65fF
C4130 BU_3VX2_2|A BU_3VX2_63|A 0.01fF
C4131 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<6> 0.01fF
C4132 LS_3VX2_7|A raven_soc_0|ser_rx 0.01fF
C4133 LOGIC0_3V_4|Q raven_soc_0|gpio_in<10> 0.08fF
C4134 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<27> 0.22fF
C4135 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<29> 0.10fF
C4136 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<9> 33.25fF
C4137 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pullup<13> 15.26fF
C4138 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pullup<6> 0.52fF
C4139 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<14> 0.62fF
C4140 BU_3VX2_27|A raven_soc_0|flash_io0_do 4.08fF
C4141 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pulldown<6> 0.02fF
C4142 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<10> 7.79fF
C4143 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<14> 0.02fF
C4144 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<8> 0.01fF
C4145 BU_3VX2_33|A raven_soc_0|flash_io0_di 1.81fF
C4146 BU_3VX2_0|Q raven_soc_0|gpio_outenb<8> 0.01fF
C4147 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<13> 3.26fF
C4148 AMUX2_3V_0|SEL LS_3VX2_17|A 0.01fF
C4149 raven_soc_0|gpio_pulldown<14> BU_3VX2_25|Q 0.01fF
C4150 raven_soc_0|gpio_pulldown<11> BU_3VX2_23|Q 0.01fF
C4151 raven_padframe_0|BBCUD4F_2|VDDR raven_padframe_0|BBCUD4F_2|GNDR 0.68fF
C4152 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<11> 28.51fF
C4153 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<12> 4.53fF
C4154 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<1> 2.03fF
C4155 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<0> 1.52fF
C4156 BU_3VX2_68|Q BU_3VX2_64|Q 2.98fF
C4157 VDD3V3 LS_3VX2_21|Q 0.19fF
C4158 LS_3VX2_20|A BU_3VX2_48|Q 26.24fF
C4159 VDD raven_padframe_0|FILLER20F_3|VDDR 0.71fF
C4160 BU_3VX2_20|A BU_3VX2_16|A 5.01fF
C4161 raven_padframe_0|CORNERESDF_2|VDDR raven_padframe_0|CORNERESDF_2|GNDR 0.68fF
C4162 BU_3VX2_20|A BU_3VX2_29|A 2.35fF
C4163 raven_padframe_0|APR00DF_0|VDDR adc_low 0.01fF
C4164 raven_padframe_0|APR00DF_3|VDDR raven_padframe_0|APR00DF_3|GNDO 0.13fF
C4165 raven_spi_0|CSB raven_padframe_0|ICFC_1|PO 0.04fF
C4166 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<11> 0.01fF
C4167 LS_3VX2_12|A LS_3VX2_21|A 6.53fF
C4168 LS_3VX2_2|A VDD3V3 0.45fF
C4169 raven_soc_0|ram_rdata<26> vdd 0.76fF
C4170 raven_soc_0|ext_clk BU_3VX2_52|Q 0.97fF
C4171 raven_soc_0|irq_pin apllc03_1v8_0|CLK 2.03fF
C4172 raven_soc_0|ram_wdata<13> vdd 0.90fF
C4173 BU_3VX2_52|A BU_3VX2_52|Q 0.10fF
C4174 VDD raven_padframe_0|BBCUD4F_15|VDDR 0.71fF
C4175 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<15> 0.01fF
C4176 BU_3VX2_23|A BU_3VX2_17|A 3.67fF
C4177 raven_padframe_0|FILLER20F_3|VDDR LOGIC0_3V_4|Q 0.01fF
C4178 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<9> 0.16fF
C4179 LS_3VX2_3|Q raven_soc_0|flash_csb 0.01fF
C4180 raven_spi_0|sdo_enb raven_soc_0|gpio_pulldown<15> 1.15fF
C4181 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<11> 0.01fF
C4182 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<11> 21.09fF
C4183 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<15> 0.86fF
C4184 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<12> 0.67fF
C4185 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<14> 0.40fF
C4186 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<6> 0.01fF
C4187 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<7> 0.01fF
C4188 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<13> 0.02fF
C4189 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<12> 5.82fF
C4190 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<9> 0.01fF
C4191 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<5> 0.01fF
C4192 BU_3VX2_7|A VDD3V3 0.21fF
C4193 BU_3VX2_6|A BU_3VX2_5|Q 0.16fF
C4194 BU_3VX2_38|A BU_3VX2_35|Q 0.16fF
C4195 LS_3VX2_24|A LS_3VX2_20|A 11.21fF
C4196 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<10> 0.01fF
C4197 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<14> 4.32fF
C4198 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<29> 3.45fF
C4199 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<6> 0.33fF
C4200 BU_3VX2_13|Q BU_3VX2_32|Q 0.20fF
C4201 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<24> 19.98fF
C4202 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<3> 32.49fF
C4203 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<31> 1.27fF
C4204 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<2> 8.01fF
C4205 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<13> 1.29fF
C4206 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io1_di 22.32fF
C4207 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<4> 8.58fF
C4208 BU_3VX2_6|Q BU_3VX2_4|Q 25.25fF
C4209 raven_soc_0|flash_io3_do raven_soc_0|flash_io0_di 54.08fF
C4210 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<17> 29.79fF
C4211 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<2> 2.51fF
C4212 BU_3VX2_21|Q BU_3VX2_70|Q 2.80fF
C4213 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<21> 55.00fF
C4214 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<22> 0.02fF
C4215 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<18> 0.01fF
C4216 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<25> 0.01fF
C4217 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<19> 0.01fF
C4218 raven_soc_0|flash_io2_do raven_soc_0|flash_io0_oeb 36.78fF
C4219 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<26> 0.01fF
C4220 BU_3VX2_4|Q BU_3VX2_7|Q 16.68fF
C4221 BU_3VX2_70|Q BU_3VX2_8|Q 1.06fF
C4222 BU_3VX2_11|Q BU_3VX2_22|Q 3.97fF
C4223 BU_3VX2_36|Q BU_3VX2_33|Q 0.76fF
C4224 LS_3VX2_17|A BU_3VX2_61|Q 25.89fF
C4225 BU_3VX2_28|Q BU_3VX2_27|Q 215.61fF
C4226 BU_3VX2_72|Q apllc03_1v8_0|B_CP 8.05fF
C4227 raven_padframe_0|BBCUD4F_15|VDDR LOGIC0_3V_4|Q 0.01fF
C4228 LOGIC0_3V_4|Q raven_soc_0|gpio_in<0> 0.09fF
C4229 raven_padframe_0|BBCUD4F_12|GNDR raven_padframe_0|BBCUD4F_12|GNDO 0.81fF
C4230 LOGIC0_3V_4|Q raven_soc_0|flash_csb 0.27fF
C4231 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<5> 0.01fF
C4232 raven_spi_0|SDO raven_soc_0|flash_io3_oeb 0.46fF
C4233 BU_3VX2_6|A raven_soc_0|flash_io1_di 0.03fF
C4234 raven_padframe_0|FILLER50F_2|VDDR raven_padframe_0|FILLER50F_2|GNDR 0.68fF
C4235 LS_3VX2_5|Q LS_3VX2_22|A 0.01fF
C4236 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<7> 0.01fF
C4237 adc_low BU_3VX2_52|A 0.06fF
C4238 VDD raven_padframe_0|aregc01_3v3_0|m4_92500_31172# 0.12fF
C4239 VDD raven_padframe_0|FILLER20F_4|GNDO 0.07fF
C4240 raven_soc_0|gpio_pulldown<10> BU_3VX2_25|Q 0.01fF
C4241 raven_soc_0|gpio_pulldown<12> BU_3VX2_27|Q 0.01fF
C4242 AMUX4_3V_0|AIN1 vdd 1.04fF
C4243 BU_3VX2_16|A BU_3VX2_14|Q 0.03fF
C4244 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<8> 0.58fF
C4245 BU_3VX2_63|Q raven_soc_0|flash_io3_do 0.17fF
C4246 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<6> 1.34fF
C4247 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<15> 321.82fF
C4248 LS_3VX2_24|Q vdd 1.20fF
C4249 raven_soc_0|gpio_outenb<2> BU_3VX2_24|Q 0.01fF
C4250 BU_3VX2_44|A BU_3VX2_43|A 4.81fF
C4251 raven_padframe_0|BT4F_1|GNDR raven_padframe_0|BT4F_1|VDDO 0.09fF
C4252 BU_3VX2_20|A LS_3VX2_3|Q 0.01fF
C4253 BU_3VX2_23|A BU_3VX2_12|A 1.90fF
C4254 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<9> 0.16fF
C4255 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<10> 0.01fF
C4256 raven_padframe_0|BBCUD4F_1|GNDR raven_padframe_0|BBCUD4F_1|VDDO 0.09fF
C4257 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<13> 0.01fF
C4258 BU_3VX2_63|Q raven_soc_0|gpio_out<14> 0.01fF
C4259 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<10> 7.31fF
C4260 raven_soc_0|flash_csb raven_soc_0|flash_io1_oeb 83.48fF
C4261 LOGIC0_3V_0|Q LOGIC1_3V_3|Q 0.01fF
C4262 BU_3VX2_19|Q vdd 1.22fF
C4263 BU_3VX2_35|Q BU_3VX2_23|Q 0.01fF
C4264 BU_3VX2_18|Q vdd 0.79fF
C4265 BU_3VX2_31|Q BU_3VX2_26|Q 9.50fF
C4266 BU_3VX2_64|Q BU_3VX2_24|Q 0.02fF
C4267 LS_3VX2_16|A BU_3VX2_57|Q 13.97fF
C4268 BU_3VX2_5|Q BU_3VX2_25|Q 0.02fF
C4269 AMUX4_3V_4|AIN2 BU_3VX2_54|Q 0.01fF
C4270 AMUX4_3V_3|SEL[0] apllc03_1v8_0|CLK 23.51fF
C4271 LS_3VX2_7|Q LS_3VX2_11|Q 13.67fF
C4272 BU_3VX2_17|A IN_3VX2_1|A 1.63fF
C4273 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<8> 0.58fF
C4274 raven_soc_0|ram_wdata<19> raven_soc_0|ram_rdata<16> 0.02fF
C4275 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<0> 8.44fF
C4276 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<16> 12.37fF
C4277 raven_soc_0|ram_wdata<29> raven_soc_0|ram_rdata<13> 0.02fF
C4278 BU_3VX2_46|A BU_3VX2_42|A 0.24fF
C4279 BU_3VX2_45|A LS_3VX2_27|Q 0.23fF
C4280 BU_3VX2_50|A BU_3VX2_50|Q 0.10fF
C4281 BU_3VX2_57|A BU_3VX2_59|Q 0.04fF
C4282 AMUX4_3V_1|SEL[0] LS_3VX2_15|A 8.87fF
C4283 raven_soc_0|flash_io1_di BU_3VX2_25|Q 0.01fF
C4284 raven_soc_0|flash_io2_oeb BU_3VX2_28|Q 0.01fF
C4285 LS_3VX2_15|Q BU_3VX2_60|Q 0.63fF
C4286 raven_soc_0|flash_io3_oeb BU_3VX2_26|Q 0.01fF
C4287 raven_soc_0|flash_io2_do BU_3VX2_29|Q 0.01fF
C4288 BU_3VX2_47|Q BU_3VX2_48|Q 221.49fF
C4289 raven_padframe_0|FILLER01F_0|VDDR raven_padframe_0|FILLER01F_0|GNDO 0.13fF
C4290 raven_padframe_0|aregc01_3v3_1|m4_92500_28769# raven_padframe_0|aregc01_3v3_1|GNDO 0.04fF
C4291 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<8> 0.01fF
C4292 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<5> 0.98fF
C4293 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<13> 8.48fF
C4294 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<9> 30.80fF
C4295 BU_3VX2_10|A raven_soc_0|flash_io2_oeb 0.01fF
C4296 LS_3VX2_9|A VDD3V3 0.51fF
C4297 LS_3VX2_12|Q LS_3VX2_19|A 0.01fF
C4298 LS_3VX2_6|Q vdd 0.13fF
C4299 VDD raven_padframe_0|APR00DF_5|VDDR 0.71fF
C4300 LS_3VX2_7|A BU_3VX2_72|Q 0.89fF
C4301 VDD raven_padframe_0|BBCUD4F_13|GNDR 0.16fF
C4302 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<5> 0.64fF
C4303 raven_soc_0|gpio_pullup<12> BU_3VX2_40|Q 0.02fF
C4304 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<10> 0.01fF
C4305 BU_3VX2_0|Q raven_soc_0|gpio_in<15> 0.01fF
C4306 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<14> 0.02fF
C4307 raven_soc_0|gpio_pullup<11> raven_soc_0|ext_clk 0.01fF
C4308 raven_soc_0|gpio_pullup<15> VDD3V3 2.66fF
C4309 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<28> 2.31fF
C4310 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<0> 0.63fF
C4311 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<19> 2.43fF
C4312 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<11> 16.65fF
C4313 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<20> 136.22fF
C4314 LS_3VX2_21|A BU_3VX2_46|Q 10.04fF
C4315 BU_3VX2_10|A BU_3VX2_6|A 3.34fF
C4316 BU_3VX2_20|A raven_soc_0|flash_io1_oeb 0.01fF
C4317 BU_3VX2_8|A raven_soc_0|flash_io0_di 0.01fF
C4318 AMUX4_3V_4|AOUT AMUX4_3V_4|AIN2 1.05fF
C4319 BU_3VX2_5|A raven_soc_0|flash_io3_do 0.03fF
C4320 BU_3VX2_0|A raven_soc_0|flash_io2_oeb 4.11fF
C4321 LS_3VX2_8|Q vdd 0.08fF
C4322 LOGIC0_3V_4|Q raven_soc_0|gpio_in<13> 0.08fF
C4323 IN_3VX2_1|A raven_soc_0|gpio_pulldown<7> 0.01fF
C4324 BU_3VX2_31|A raven_soc_0|flash_io2_di 4.02fF
C4325 raven_spi_0|sdo_enb raven_soc_0|flash_io3_di 1.22fF
C4326 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<6> 9.46fF
C4327 LS_3VX2_24|A BU_3VX2_47|Q 5.67fF
C4328 BU_3VX2_27|A raven_soc_0|flash_io1_di 0.01fF
C4329 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pulldown<6> 0.02fF
C4330 LS_3VX2_3|A BU_3VX2_71|Q 120.71fF
C4331 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<12> 3.71fF
C4332 raven_padframe_0|FILLER20F_3|VDDR raven_padframe_0|FILLER20F_3|GNDR 0.68fF
C4333 raven_padframe_0|BBCUD4F_0|VDDR raven_padframe_0|BBCUD4F_0|GNDO 0.13fF
C4334 BU_3VX2_6|A BU_3VX2_0|A 0.05fF
C4335 LS_3VX2_12|Q adc_low 0.12fF
C4336 IN_3VX2_1|A BU_3VX2_12|A 0.01fF
C4337 LS_3VX2_12|A LS_3VX2_27|A 7.46fF
C4338 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<14> 2.65fF
C4339 LOGIC0_3V_1|Q raven_spi_0|SDI 2.16fF
C4340 raven_soc_0|ram_wdata<12> vdd 0.75fF
C4341 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<9> 0.01fF
C4342 raven_soc_0|gpio_pulldown<1> BU_3VX2_63|Q 0.13fF
C4343 BU_3VX2_31|A raven_soc_0|gpio_pulldown<11> 0.01fF
C4344 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<13> 0.01fF
C4345 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<6> 0.05fF
C4346 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<10> 9.30fF
C4347 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<7> 0.02fF
C4348 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<14> 0.02fF
C4349 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<11> 50.22fF
C4350 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<12> 5.60fF
C4351 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<11> 0.02fF
C4352 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<12> 5.28fF
C4353 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<15> 0.02fF
C4354 BU_3VX2_0|Q raven_soc_0|gpio_out<13> 0.01fF
C4355 raven_soc_0|gpio_out<1> BU_3VX2_29|Q 0.01fF
C4356 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<8> 3.46fF
C4357 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<9> 0.15fF
C4358 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<6> 0.17fF
C4359 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<22> 1.05fF
C4360 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<20> 51.13fF
C4361 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<24> 61.07fF
C4362 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<5> 0.01fF
C4363 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<23> 1.86fF
C4364 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<31> 0.08fF
C4365 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<18> 8.28fF
C4366 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<6> 8.12fF
C4367 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<3> 0.01fF
C4368 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<2> 0.28fF
C4369 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<25> 4.68fF
C4370 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<2> 1.60fF
C4371 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<1> 0.03fF
C4372 BU_3VX2_6|Q BU_3VX2_3|Q 19.34fF
C4373 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<19> 0.05fF
C4374 BU_3VX2_19|Q BU_3VX2_70|Q 0.01fF
C4375 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<12> 1.37fF
C4376 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<14> 6.07fF
C4377 BU_3VX2_35|Q BU_3VX2_4|Q 5.78fF
C4378 BU_3VX2_12|Q BU_3VX2_37|Q 3.05fF
C4379 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<8> 3.20fF
C4380 BU_3VX2_70|Q BU_3VX2_18|Q 3.36fF
C4381 BU_3VX2_3|Q BU_3VX2_7|Q 10.23fF
C4382 AMUX4_3V_4|SEL[0] AMUX4_3V_4|SEL[1] 163.70fF
C4383 BU_3VX2_14|Q BU_3VX2_67|Q 16.36fF
C4384 AMUX4_3V_1|SEL[0] AMUX4_3V_1|SEL[1] 195.58fF
C4385 BU_3VX2_32|Q BU_3VX2_69|Q 0.49fF
C4386 LS_3VX2_17|A LS_3VX2_15|A 36.64fF
C4387 BU_3VX2_25|Q BU_3VX2_28|Q 77.00fF
C4388 vdd BU_3VX2_27|Q 1.62fF
C4389 BU_3VX2_24|Q apllc03_1v8_0|B_VCO 0.76fF
C4390 BU_3VX2_26|Q apllc03_1v8_0|CLK 7.85fF
C4391 raven_spi_0|CSB LOGIC0_3V_3|Q 1.49fF
C4392 BU_3VX2_25|A BU_3VX2_17|A 2.70fF
C4393 raven_padframe_0|CORNERESDF_0|VDDR raven_padframe_0|CORNERESDF_0|GNDO 0.13fF
C4394 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<1> 9.58fF
C4395 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<14> 0.01fF
C4396 BU_3VX2_32|A vdd 0.16fF
C4397 LS_3VX2_14|A AMUX4_3V_4|AIN2 1.38fF
C4398 LS_3VX2_7|A AMUX4_3V_1|SEL[0] 10.60fF
C4399 raven_soc_0|gpio_pulldown<12> BU_3VX2_25|Q 0.01fF
C4400 raven_soc_0|ram_rdata<11> raven_soc_0|ram_addr<0> 0.01fF
C4401 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<1> 0.09fF
C4402 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<15> 3.80fF
C4403 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<17> 27.00fF
C4404 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<31> 0.02fF
C4405 BU_3VX2_71|Q raven_soc_0|flash_io1_do 0.05fF
C4406 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<14> 22.20fF
C4407 raven_soc_0|gpio_out<3> VDD3V3 0.45fF
C4408 raven_soc_0|gpio_pulldown<8> raven_soc_0|ext_clk 0.01fF
C4409 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<7> 0.01fF
C4410 BU_3VX2_27|A BU_3VX2_28|Q 0.03fF
C4411 raven_soc_0|gpio_in<2> BU_3VX2_27|Q 0.01fF
C4412 AMUX2_3V_0|SEL BU_3VX2_42|Q 9.20fF
C4413 adc_high BU_3VX2_59|Q 0.07fF
C4414 VDD raven_padframe_0|GNDORPADF_3|VDDR 0.71fF
C4415 BU_3VX2_10|A BU_3VX2_27|A 0.01fF
C4416 LS_3VX2_14|Q LS_3VX2_4|A 0.54fF
C4417 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<4> 0.70fF
C4418 raven_soc_0|gpio_outenb<3> LS_3VX2_3|A 0.01fF
C4419 BU_3VX2_22|A raven_soc_0|flash_io2_di 0.01fF
C4420 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<4> 1.84fF
C4421 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<13> 0.22fF
C4422 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<6> 0.01fF
C4423 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<8> 0.01fF
C4424 raven_soc_0|gpio_in<15> raven_soc_0|irq_pin 0.01fF
C4425 raven_soc_0|irq_pin BU_3VX2_43|Q 24.50fF
C4426 AMUX4_3V_4|AIN2 BU_3VX2_56|Q 0.01fF
C4427 AMUX4_3V_4|SEL[1] vdd 5.98fF
C4428 BU_3VX2_8|A BU_3VX2_5|A 5.00fF
C4429 raven_padframe_0|GNDORPADF_3|VDDR LOGIC0_3V_4|Q 0.01fF
C4430 raven_padframe_0|ICFC_1|VDD3 LOGIC0_3V_4|Q 0.04fF
C4431 LS_3VX2_11|Q LS_3VX2_4|Q 0.75fF
C4432 BU_3VX2_25|A BU_3VX2_12|A 1.59fF
C4433 BU_3VX2_0|A BU_3VX2_27|A 0.01fF
C4434 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<1> 0.01fF
C4435 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_out<2> 37.64fF
C4436 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<10> 0.01fF
C4437 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<13> 0.21fF
C4438 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<29> 0.01fF
C4439 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<9> 21.03fF
C4440 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<16> 0.01fF
C4441 raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<27> 61.91fF
C4442 raven_soc_0|ram_wdata<17> raven_soc_0|ram_rdata<17> 0.48fF
C4443 raven_soc_0|ram_rdata<2> raven_soc_0|ram_addr<0> 1.03fF
C4444 raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<31> 8.49fF
C4445 LS_3VX2_15|Q BU_3VX2_62|Q 5.34fF
C4446 raven_soc_0|flash_io2_oeb vdd 3.49fF
C4447 AMUX4_3V_1|SEL[1] LS_3VX2_17|A 0.43fF
C4448 BU_3VX2_50|A LS_3VX2_27|Q 0.10fF
C4449 BU_3VX2_49|A LS_3VX2_20|Q 0.17fF
C4450 BU_3VX2_48|A BU_3VX2_43|A 0.38fF
C4451 raven_soc_0|flash_io3_do BU_3VX2_24|Q 0.01fF
C4452 raven_soc_0|gpio_in<11> BU_3VX2_27|Q 0.01fF
C4453 BU_3VX2_50|A BU_3VX2_48|Q 0.04fF
C4454 AMUX4_3V_3|AOUT AMUX4_3V_4|AOUT 41.20fF
C4455 BU_3VX2_35|A BU_3VX2_71|A 0.01fF
C4456 aopac01_3v3_0|IB acsoc02_3v3_0|CS_8U 0.25fF
C4457 raven_soc_0|gpio_out<0> BU_3VX2_63|Q 0.01fF
C4458 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<7> 0.01fF
C4459 raven_padframe_0|axtoc02_3v3_0|m4_55000_31172# raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# 0.02fF
C4460 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<6> 0.01fF
C4461 BU_3VX2_63|Q raven_soc_0|gpio_out<12> 0.01fF
C4462 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<10> 6.74fF
C4463 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<15> 113.97fF
C4464 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<6> 0.01fF
C4465 BU_3VX2_7|A BU_3VX2_8|Q 0.03fF
C4466 BU_3VX2_6|A vdd 0.13fF
C4467 BU_3VX2_18|A BU_3VX2_16|Q 0.03fF
C4468 LS_3VX2_12|Q LS_3VX2_22|A 0.01fF
C4469 LS_3VX2_7|A LS_3VX2_17|A 0.01fF
C4470 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<13> 197.40fF
C4471 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<12> 0.02fF
C4472 raven_soc_0|gpio_outenb<0> BU_3VX2_40|Q 0.02fF
C4473 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<7> 0.01fF
C4474 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<5> 0.01fF
C4475 BU_3VX2_0|Q raven_soc_0|gpio_in<14> 0.01fF
C4476 raven_soc_0|gpio_outenb<9> BU_3VX2_27|Q 0.01fF
C4477 raven_soc_0|gpio_outenb<13> apllc03_1v8_0|CLK 0.01fF
C4478 raven_soc_0|gpio_out<14> BU_3VX2_24|Q 0.01fF
C4479 BU_3VX2_4|Q BU_3VX2_23|Q 0.37fF
C4480 BU_3VX2_32|Q BU_3VX2_29|Q 5.49fF
C4481 BU_3VX2_70|Q BU_3VX2_27|Q 0.40fF
C4482 LS_3VX2_27|A BU_3VX2_46|Q 10.18fF
C4483 BU_3VX2_11|Q apllc03_1v8_0|CLK 0.01fF
C4484 raven_spi_0|CSB VDD3V3 0.19fF
C4485 BU_3VX2_18|A raven_soc_0|flash_io3_di 0.01fF
C4486 BU_3VX2_40|A raven_soc_0|flash_io2_oeb 0.01fF
C4487 raven_padframe_0|BBC4F_3|VDDR raven_padframe_0|BBC4F_3|GNDR 0.68fF
C4488 BU_3VX2_13|A raven_soc_0|flash_io3_do 0.01fF
C4489 raven_soc_0|gpio_in<2> raven_soc_0|flash_io2_oeb 16.20fF
C4490 LS_3VX2_8|A BU_3VX2_51|Q 5.04fF
C4491 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pulldown<6> 1.87fF
C4492 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<5> 5.69fF
C4493 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<0> 38.64fF
C4494 BU_3VX2_0|Q raven_soc_0|gpio_pullup<6> 0.07fF
C4495 LS_3VX2_3|A raven_soc_0|gpio_pullup<14> 0.33fF
C4496 BU_3VX2_33|A raven_soc_0|gpio_out<15> 11.14fF
C4497 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pulldown<7> 0.01fF
C4498 raven_padframe_0|FILLER02F_0|VDDR raven_padframe_0|FILLER02F_0|GNDR 0.68fF
C4499 BU_3VX2_41|A BU_3VX2_45|A 2.55fF
C4500 BU_3VX2_41|A BU_3VX2_47|Q 0.03fF
C4501 BU_3VX2_7|A BU_3VX2_19|A 0.95fF
C4502 BU_3VX2_6|A BU_3VX2_40|A 0.79fF
C4503 raven_spi_0|SDO raven_spi_0|sdo_enb 139.07fF
C4504 BU_3VX2_38|A BU_3VX2_31|A 0.01fF
C4505 LS_3VX2_5|Q LS_3VX2_5|A 0.05fF
C4506 BU_3VX2_23|A raven_soc_0|flash_clk 3.73fF
C4507 BU_3VX2_70|A BU_3VX2_36|A 1.56fF
C4508 BU_3VX2_21|A raven_soc_0|flash_io2_di 0.12fF
C4509 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<3> 0.01fF
C4510 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<6> 0.01fF
C4511 raven_soc_0|gpio_in<4> raven_soc_0|flash_io1_di 0.19fF
C4512 IN_3VX2_1|A BU_3VX2_59|Q 0.01fF
C4513 raven_soc_0|gpio_out<11> BU_3VX2_29|Q 0.01fF
C4514 BU_3VX2_53|A BU_3VX2_55|Q 0.04fF
C4515 raven_soc_0|irq_pin BU_3VX2_50|Q 7.30fF
C4516 raven_soc_0|irq_pin raven_padframe_0|ICF_1|PO 0.04fF
C4517 BU_3VX2_23|A BU_3VX2_9|A 0.01fF
C4518 BU_3VX2_68|A BU_3VX2_67|A 24.99fF
C4519 BU_3VX2_4|A BU_3VX2_17|A 0.78fF
C4520 LS_3VX2_7|Q LS_3VX2_8|A 0.16fF
C4521 LOGIC1_3V_2|Q LOGIC0_3V_3|Q 2.89fF
C4522 BU_3VX2_0|A BU_3VX2_64|A 2.79fF
C4523 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<12> 1.19fF
C4524 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<7> 0.01fF
C4525 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<11> 23.43fF
C4526 BU_3VX2_0|Q raven_soc_0|gpio_outenb<15> 0.01fF
C4527 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<11> 0.01fF
C4528 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<15> 0.02fF
C4529 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<7> 0.01fF
C4530 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<12> 5.11fF
C4531 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<24> 0.37fF
C4532 AMUX4_3V_3|SEL[1] BU_3VX2_66|Q 4.24fF
C4533 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<21> 0.40fF
C4534 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<22> 0.46fF
C4535 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<30> 0.19fF
C4536 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<14> 0.21fF
C4537 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<23> 3.71fF
C4538 BU_3VX2_14|Q BU_3VX2_65|Q 19.72fF
C4539 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<12> 9.45fF
C4540 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<25> 0.81fF
C4541 BU_3VX2_37|Q BU_3VX2_5|Q 12.30fF
C4542 raven_soc_0|gpio_in<1> LOGIC0_3V_4|Q 0.09fF
C4543 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<1> 0.06fF
C4544 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<15> 0.19fF
C4545 raven_soc_0|gpio_out<15> raven_soc_0|flash_io3_do 1.99fF
C4546 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<8> 0.01fF
C4547 BU_3VX2_35|Q BU_3VX2_3|Q 7.56fF
C4548 BU_3VX2_40|Q raven_soc_0|flash_io0_do 0.01fF
C4549 vdd BU_3VX2_25|Q 0.69fF
C4550 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<2> 8.09fF
C4551 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<5> 0.01fF
C4552 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<2> 3.41fF
C4553 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_out<9> 0.22fF
C4554 raven_spi_0|SDO raven_soc_0|gpio_in<15> 1.54fF
C4555 AMUX4_3V_1|AIN1 BU_3VX2_58|A 0.02fF
C4556 BU_3VX2_12|A BU_3VX2_13|Q 0.03fF
C4557 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<23> 0.08fF
C4558 BU_3VX2_71|Q raven_soc_0|gpio_in<10> 0.21fF
C4559 raven_soc_0|gpio_out<14> raven_soc_0|gpio_out<15> 32.02fF
C4560 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<19> 0.01fF
C4561 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<20> 0.01fF
C4562 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<22> 0.02fF
C4563 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<29> 0.02fF
C4564 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<25> 2.00fF
C4565 AMUX4_3V_0|AIN1 LS_3VX2_21|Q 1.14fF
C4566 IN_3VX2_1|Q AMUX4_3V_1|SEL[0] 0.01fF
C4567 BU_3VX2_15|A BU_3VX2_12|Q 0.02fF
C4568 LS_3VX2_9|Q VDD3V3 0.21fF
C4569 LS_3VX2_14|Q vdd 0.96fF
C4570 VDD raven_padframe_0|FILLER01F_0|VDDR 0.71fF
C4571 BU_3VX2_26|A raven_soc_0|flash_io3_oeb 2.91fF
C4572 raven_soc_0|gpio_pulldown<14> BU_3VX2_40|Q 0.03fF
C4573 BU_3VX2_63|Q raven_soc_0|gpio_pullup<5> 0.04fF
C4574 raven_soc_0|gpio_in<2> BU_3VX2_25|Q 0.01fF
C4575 BU_3VX2_31|A BU_3VX2_23|Q 73.50fF
C4576 adc_high BU_3VX2_61|Q 0.06fF
C4577 raven_soc_0|gpio_pulldown<1> BU_3VX2_24|Q 0.01fF
C4578 BU_3VX2_27|A vdd 0.06fF
C4579 LS_3VX2_13|A LS_3VX2_20|A 6.43fF
C4580 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_outenb<8> 1.66fF
C4581 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<10> 0.08fF
C4582 raven_soc_0|gpio_in<5> raven_soc_0|gpio_out<14> 1.76fF
C4583 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<31> 0.47fF
C4584 raven_padframe_0|FILLER10F_1|GNDR raven_padframe_0|FILLER10F_1|VDDO 0.09fF
C4585 BU_3VX2_63|A BU_3VX2_18|A 0.01fF
C4586 BU_3VX2_2|A BU_3VX2_26|A 1.18fF
C4587 BU_3VX2_4|A BU_3VX2_12|A 1.29fF
C4588 AMUX4_3V_3|AOUT raven_soc_0|flash_io0_oeb 4.79fF
C4589 BU_3VX2_3|A raven_soc_0|flash_io0_do 0.01fF
C4590 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<13> 0.01fF
C4591 BU_3VX2_71|A raven_soc_0|flash_io3_di 0.01fF
C4592 raven_soc_0|gpio_pullup<2> BU_3VX2_27|Q 0.01fF
C4593 BU_3VX2_15|A raven_soc_0|flash_io0_do 0.01fF
C4594 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<13> 0.27fF
C4595 IN_3VX2_1|A raven_soc_0|flash_clk 40.55fF
C4596 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<6> 0.83fF
C4597 BU_3VX2_11|A raven_soc_0|flash_io3_oeb 0.01fF
C4598 raven_soc_0|gpio_in<14> raven_soc_0|irq_pin 0.01fF
C4599 raven_padframe_0|ICFC_2|VDDR raven_padframe_0|ICFC_2|VDD3 0.71fF
C4600 BU_3VX2_23|A BU_3VX2_28|A 7.89fF
C4601 BU_3VX2_8|A BU_3VX2_13|A 2.47fF
C4602 BU_3VX2_9|A IN_3VX2_1|A 0.01fF
C4603 BU_3VX2_2|A LOGIC0_3V_3|Q 0.28fF
C4604 LS_3VX2_10|A LS_3VX2_6|A 155.16fF
C4605 BU_3VX2_0|A BU_3VX2_66|A 0.95fF
C4606 BU_3VX2_2|A BU_3VX2_11|A 1.75fF
C4607 BU_3VX2_40|A BU_3VX2_27|A 0.13fF
C4608 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<12> 0.01fF
C4609 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<1> 24.87fF
C4610 raven_soc_0|gpio_in<0> BU_3VX2_71|Q 0.02fF
C4611 raven_soc_0|flash_csb BU_3VX2_71|Q 0.01fF
C4612 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<31> 6.52fF
C4613 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<7> 5.07fF
C4614 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<27> 0.01fF
C4615 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<21> 0.01fF
C4616 BU_3VX2_24|A BU_3VX2_35|A 0.01fF
C4617 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<17> 0.01fF
C4618 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<0> 0.01fF
C4619 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<25> 0.01fF
C4620 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<17> 0.01fF
C4621 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<13> 3.90fF
C4622 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<16> 12.32fF
C4623 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<21> 59.11fF
C4624 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<25> 180.29fF
C4625 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<22> 16.58fF
C4626 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<29> 4.71fF
C4627 raven_soc_0|ram_wdata<15> raven_soc_0|ram_rdata<1> 0.02fF
C4628 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<31> 0.01fF
C4629 LS_3VX2_19|A BU_3VX2_55|Q 7.81fF
C4630 raven_soc_0|gpio_in<8> apllc03_1v8_0|CLK 0.02fF
C4631 LS_3VX2_16|Q LS_3VX2_16|A 0.06fF
C4632 raven_soc_0|gpio_in<15> BU_3VX2_26|Q 0.01fF
C4633 raven_soc_0|gpio_in<11> BU_3VX2_25|Q 0.01fF
C4634 raven_soc_0|gpio_in<12> BU_3VX2_29|Q 0.01fF
C4635 raven_soc_0|gpio_in<7> BU_3VX2_28|Q 0.01fF
C4636 BU_3VX2_55|Q BU_3VX2_52|Q 50.22fF
C4637 AMUX4_3V_0|SEL[1] BU_3VX2_44|Q 58.76fF
C4638 BU_3VX2_44|Q BU_3VX2_51|Q 15.10fF
C4639 LS_3VX2_20|Q BU_3VX2_46|Q 0.11fF
C4640 raven_padframe_0|VDDPADFC_0|GNDR raven_padframe_0|VDDPADFC_0|VDDO 0.09fF
C4641 LOGIC1_3V_1|Q LOGIC0_3V_4|Q 0.17fF
C4642 raven_padframe_0|aregc01_3v3_1|m4_92500_29333# raven_padframe_0|aregc01_3v3_1|m4_92500_29057# 0.11fF
C4643 raven_padframe_0|aregc01_3v3_1|m4_92500_30133# raven_padframe_0|aregc01_3v3_1|m4_92500_28769# 0.01fF
C4644 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<11> 53.61fF
C4645 BU_3VX2_63|Q raven_soc_0|gpio_outenb<12> 0.01fF
C4646 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<8> 0.01fF
C4647 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<10> 5.13fF
C4648 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<7> 0.01fF
C4649 LOGIC1_3V_2|Q VDD3V3 0.06fF
C4650 raven_soc_0|gpio_pulldown<10> BU_3VX2_40|Q 0.04fF
C4651 LS_3VX2_3|A raven_soc_0|gpio_in<9> 0.01fF
C4652 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<7> 0.01fF
C4653 BU_3VX2_37|Q BU_3VX2_28|Q 0.37fF
C4654 BU_3VX2_3|Q BU_3VX2_23|Q 0.45fF
C4655 raven_soc_0|gpio_pullup<13> apllc03_1v8_0|CLK 0.01fF
C4656 raven_soc_0|gpio_outenb<9> BU_3VX2_25|Q 0.01fF
C4657 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<4> 7.35fF
C4658 IN_3VX2_1|Q LS_3VX2_17|A 0.01fF
C4659 raven_padframe_0|BBC4F_1|VDDR raven_padframe_0|BBC4F_1|GNDO 0.13fF
C4660 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<8> 0.73fF
C4661 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<7> 3.44fF
C4662 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<3> 0.57fF
C4663 BU_3VX2_0|Q AMUX4_3V_3|SEL[1] 11.17fF
C4664 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<5> 0.01fF
C4665 adc_low BU_3VX2_55|Q 0.05fF
C4666 raven_soc_0|gpio_outenb<2> raven_soc_0|ext_clk 0.01fF
C4667 BU_3VX2_64|A vdd 0.22fF
C4668 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<19> 8.26fF
C4669 BU_3VX2_51|A BU_3VX2_46|A 0.69fF
C4670 BU_3VX2_49|A BU_3VX2_47|A 3.67fF
C4671 BU_3VX2_50|A BU_3VX2_41|A 1.23fF
C4672 raven_padframe_0|APR00DF_4|VDDO raven_padframe_0|APR00DF_4|GNDO 2.28fF
C4673 LS_3VX2_12|A BU_3VX2_53|Q 10.91fF
C4674 BU_3VX2_22|A BU_3VX2_23|Q 0.03fF
C4675 raven_soc_0|gpio_out<0> BU_3VX2_24|Q 0.01fF
C4676 BU_3VX2_17|A raven_soc_0|flash_io0_oeb 0.01fF
C4677 IN_3VX2_1|A BU_3VX2_61|Q 0.01fF
C4678 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<3> 1.52fF
C4679 raven_soc_0|gpio_out<13> BU_3VX2_26|Q 0.01fF
C4680 raven_soc_0|ram_wenb vdd 0.32fF
C4681 raven_soc_0|gpio_out<5> apllc03_1v8_0|CLK 0.01fF
C4682 raven_soc_0|gpio_out<12> BU_3VX2_24|Q 0.01fF
C4683 raven_soc_0|gpio_outenb<14> BU_3VX2_27|Q 0.01fF
C4684 BU_3VX2_73|Q VDD3V3 0.08fF
C4685 raven_soc_0|irq_pin BU_3VX2_48|Q 8.90fF
C4686 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<13> 0.01fF
C4687 VDD3V3 raven_padframe_0|VDDORPADF_2|GNDO 2.41fF
C4688 BU_3VX2_63|A BU_3VX2_71|A 2.55fF
C4689 BU_3VX2_32|A BU_3VX2_69|A 0.55fF
C4690 IN_3VX2_1|A BU_3VX2_28|A 35.36fF
C4691 raven_padframe_0|axtoc02_3v3_0|XO XO 2.43fF
C4692 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<6> 0.99fF
C4693 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<4> 13.17fF
C4694 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<9> 0.15fF
C4695 BU_3VX2_25|A raven_soc_0|flash_clk 4.15fF
C4696 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<7> 0.01fF
C4697 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<12> 0.02fF
C4698 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<5> 0.01fF
C4699 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<7> 0.01fF
C4700 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<6> 0.02fF
C4701 AMUX4_3V_3|SEL[1] BU_3VX2_30|Q 0.64fF
C4702 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<12> 4.39fF
C4703 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<5> 0.27fF
C4704 AMUX4_3V_3|SEL[1] BU_3VX2_16|Q 0.18fF
C4705 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<7> 0.15fF
C4706 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<1> 0.04fF
C4707 BU_3VX2_40|Q raven_soc_0|flash_io1_di 17.56fF
C4708 raven_soc_0|ser_tx raven_soc_0|irq_pin 291.01fF
C4709 raven_soc_0|flash_io3_oeb VDD3V3 11.48fF
C4710 AMUX4_3V_0|SEL[1] vdd 4.74fF
C4711 BU_3VX2_51|Q vdd 3.84fF
C4712 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<1> 40.99fF
C4713 raven_soc_0|gpio_in<12> raven_padframe_0|BBCUD4F_12|PO 0.04fF
C4714 BU_3VX2_9|A BU_3VX2_25|A 0.01fF
C4715 raven_padframe_0|FILLER20F_8|GNDR raven_padframe_0|FILLER20F_8|VDDO 0.09fF
C4716 raven_padframe_0|VDDPADF_1|VDDR LOGIC0_3V_4|Q 0.01fF
C4717 BU_3VX2_23|A BU_3VX2_14|A 2.25fF
C4718 raven_spi_0|SDI LOGIC0_3V_2|Q 1.58fF
C4719 BU_3VX2_35|A BU_3VX2_29|A 0.01fF
C4720 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_in<0> 0.01fF
C4721 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<7> 0.01fF
C4722 raven_padframe_0|aregc01_3v3_0|m4_0_30133# raven_padframe_0|aregc01_3v3_0|GNDR 0.07fF
C4723 raven_padframe_0|aregc01_3v3_0|m4_92500_29333# raven_padframe_0|aregc01_3v3_0|m4_92500_28769# 0.03fF
C4724 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_outenb<5> 0.01fF
C4725 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<12> 0.28fF
C4726 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<10> 0.23fF
C4727 acmpc01_3v3_0|IBN VDD3V3 0.06fF
C4728 BU_3VX2_2|A VDD3V3 0.29fF
C4729 LS_3VX2_7|A BU_3VX2_42|Q 5.84fF
C4730 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<0> 0.11fF
C4731 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<23> 1.12fF
C4732 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<15> 10.15fF
C4733 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<11> 0.01fF
C4734 BU_3VX2_71|Q raven_soc_0|gpio_in<13> 0.51fF
C4735 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<6> 1.25fF
C4736 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<20> 11.22fF
C4737 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<8> 67.52fF
C4738 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<10> 0.01fF
C4739 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<13> 0.01fF
C4740 raven_soc_0|ram_addr<4> vdd 0.43fF
C4741 BU_3VX2_59|Q BU_3VX2_54|Q 27.77fF
C4742 BU_3VX2_58|Q BU_3VX2_55|Q 48.78fF
C4743 BU_3VX2_37|A BU_3VX2_35|A 11.11fF
C4744 LS_3VX2_7|Q vdd 0.09fF
C4745 BU_3VX2_65|A BU_3VX2_64|Q 0.16fF
C4746 BU_3VX2_12|A raven_soc_0|flash_io0_oeb 0.01fF
C4747 BU_3VX2_66|A vdd 0.22fF
C4748 raven_soc_0|gpio_outenb<4> VDD3V3 0.20fF
C4749 VDD raven_padframe_0|aregc01_3v3_1|m4_92500_31172# 0.12fF
C4750 raven_soc_0|gpio_pulldown<2> BU_3VX2_23|Q 0.09fF
C4751 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_outenb<8> 0.58fF
C4752 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<31> 0.23fF
C4753 raven_soc_0|gpio_out<10> raven_soc_0|gpio_out<14> 1.28fF
C4754 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<9> 0.87fF
C4755 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<10> 5.14fF
C4756 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<6> 0.05fF
C4757 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<24> 0.02fF
C4758 BU_3VX2_3|Q BU_3VX2_4|Q 75.09fF
C4759 BU_3VX2_14|Q BU_3VX2_36|Q 1.99fF
C4760 raven_padframe_0|BT4F_0|GNDR raven_padframe_0|BT4F_0|VDDO 0.09fF
C4761 BU_3VX2_24|A raven_soc_0|flash_io3_di 0.01fF
C4762 abgpc01_3v3_0|VBGVTN AMUX4_3V_4|AIN3 0.34fF
C4763 LS_3VX2_4|Q LS_3VX2_4|A 0.05fF
C4764 raven_soc_0|gpio_pullup<0> LS_3VX2_3|A 0.01fF
C4765 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<2> 0.86fF
C4766 BU_3VX2_3|A raven_soc_0|flash_io1_di 0.01fF
C4767 raven_padframe_0|BBC4F_0|VDDR raven_padframe_0|BBC4F_0|VDDO 0.06fF
C4768 BU_3VX2_15|A raven_soc_0|flash_io1_di 0.01fF
C4769 raven_soc_0|gpio_pullup<2> BU_3VX2_25|Q 0.01fF
C4770 raven_soc_0|gpio_in<3> raven_soc_0|flash_io3_do 0.78fF
C4771 LS_3VX2_6|A raven_soc_0|ser_tx 0.01fF
C4772 raven_soc_0|gpio_in<4> vdd 1.06fF
C4773 VDD raven_padframe_0|BBCUD4F_4|GNDO 0.07fF
C4774 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<15> 1.44fF
C4775 BU_3VX2_0|Q raven_soc_0|ram_rdata<19> 0.02fF
C4776 VDD raven_padframe_0|BBCUD4F_6|VDDR 0.71fF
C4777 raven_spi_0|SDO raven_soc_0|gpio_outenb<15> 1.66fF
C4778 LS_3VX2_24|A LS_3VX2_6|A 9.68fF
C4779 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<5> 0.27fF
C4780 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<14> 0.01fF
C4781 raven_soc_0|gpio_out<13> raven_soc_0|gpio_outenb<13> 192.08fF
C4782 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<14> 4.07fF
C4783 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<5> 0.10fF
C4784 raven_soc_0|gpio_out<5> raven_soc_0|gpio_outenb<8> 0.01fF
C4785 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<14> 0.01fF
C4786 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<1> 9.39fF
C4787 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<8> 0.01fF
C4788 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<9> 0.01fF
C4789 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<2> 1.52fF
C4790 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<26> 0.80fF
C4791 BU_3VX2_13|Q BU_3VX2_2|Q 3.99fF
C4792 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<13> 0.36fF
C4793 BU_3VX2_38|Q BU_3VX2_66|Q 0.98fF
C4794 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<25> 37.13fF
C4795 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<22> 22.20fF
C4796 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<21> 9.50fF
C4797 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<1> 0.01fF
C4798 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<25> 0.01fF
C4799 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<29> 5.52fF
C4800 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<19> 0.01fF
C4801 BU_3VX2_12|Q BU_3VX2_17|Q 7.87fF
C4802 BU_3VX2_22|Q BU_3VX2_8|Q 0.70fF
C4803 BU_3VX2_13|Q BU_3VX2_10|Q 13.75fF
C4804 BU_3VX2_21|Q BU_3VX2_22|Q 81.57fF
C4805 LS_3VX2_2|A AMUX4_3V_4|SEL[1] 5.68fF
C4806 raven_soc_0|ram_wdata<1> raven_soc_0|ram_rdata<1> 0.21fF
C4807 raven_soc_0|ram_wdata<0> raven_soc_0|ram_rdata<13> 0.01fF
C4808 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<19> 12.42fF
C4809 BU_3VX2_66|Q BU_3VX2_67|Q 21.39fF
C4810 BU_3VX2_67|Q BU_3VX2_20|Q 0.01fF
C4811 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<26> 5.07fF
C4812 LS_3VX2_22|A BU_3VX2_55|Q 0.02fF
C4813 BU_3VX2_1|Q BU_3VX2_68|Q 0.54fF
C4814 LS_3VX2_19|A BU_3VX2_57|Q 9.64fF
C4815 raven_soc_0|gpio_in<7> vdd 1.58fF
C4816 BU_3VX2_57|Q BU_3VX2_52|Q 38.16fF
C4817 AMUX4_3V_0|SEL[0] BU_3VX2_43|Q 56.29fF
C4818 BU_3VX2_61|A vdd 0.07fF
C4819 BU_3VX2_44|A BU_3VX2_45|Q 0.03fF
C4820 VDD3V3 apllc03_1v8_0|CLK 12.23fF
C4821 BU_3VX2_40|Q BU_3VX2_28|Q 2.17fF
C4822 raven_soc_0|gpio_in<14> BU_3VX2_26|Q 0.01fF
C4823 LS_3VX2_20|A BU_3VX2_72|Q 4.44fF
C4824 BU_3VX2_44|Q BU_3VX2_49|Q 20.65fF
C4825 VDD raven_padframe_0|BBCUD4F_0|VDDR 0.71fF
C4826 BU_3VX2_35|A LS_3VX2_3|Q 0.01fF
C4827 VDD raven_soc_0|gpio_pulldown<15> 0.24fF
C4828 raven_padframe_0|BBCUD4F_6|VDDR LOGIC0_3V_4|Q 0.01fF
C4829 BU_3VX2_25|A BU_3VX2_28|A 12.30fF
C4830 raven_padframe_0|aregc01_3v3_1|m4_0_29057# raven_padframe_0|aregc01_3v3_1|m4_0_28769# 0.11fF
C4831 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<2> 2.18fF
C4832 IN_3VX2_1|A BU_3VX2_14|A 0.01fF
C4833 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<6> 1.00fF
C4834 raven_padframe_0|axtoc02_3v3_0|m4_0_30653# raven_padframe_0|axtoc02_3v3_0|m4_0_29057# 0.01fF
C4835 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<11> 170.20fF
C4836 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<4> 0.65fF
C4837 BU_3VX2_63|Q raven_soc_0|gpio_pullup<12> 0.01fF
C4838 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<9> 0.01fF
C4839 BU_3VX2_70|A VDD3V3 0.02fF
C4840 raven_soc_0|gpio_pulldown<12> BU_3VX2_40|Q 0.04fF
C4841 BU_3VX2_37|Q vdd 1.35fF
C4842 LS_3VX2_12|A LS_3VX2_11|Q 0.16fF
C4843 raven_padframe_0|BBCUD4F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C4844 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<15> 56.35fF
C4845 BU_3VX2_7|A raven_soc_0|flash_io2_oeb 0.01fF
C4846 BU_3VX2_16|A BU_3VX2_16|Q 0.08fF
C4847 BU_3VX2_4|A BU_3VX2_2|Q 0.03fF
C4848 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<6> 0.69fF
C4849 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<7> 0.36fF
C4850 BU_3VX2_29|A BU_3VX2_30|Q 0.03fF
C4851 BU_3VX2_33|A raven_soc_0|ext_clk 1.53fF
C4852 adc_low BU_3VX2_57|Q 0.05fF
C4853 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<15> 8.40fF
C4854 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<16> 0.05fF
C4855 BU_3VX2_47|A BU_3VX2_46|Q 0.04fF
C4856 BU_3VX2_7|A BU_3VX2_6|A 22.49fF
C4857 BU_3VX2_23|A raven_soc_0|flash_io1_do 0.01fF
C4858 BU_3VX2_35|A BU_3VX2_38|Q 0.03fF
C4859 BU_3VX2_16|A raven_soc_0|flash_io3_di 0.07fF
C4860 BU_3VX2_4|A raven_soc_0|flash_clk 0.01fF
C4861 LS_3VX2_14|A BU_3VX2_59|Q 0.03fF
C4862 BU_3VX2_17|A raven_soc_0|flash_io2_do 0.01fF
C4863 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<11> 34.50fF
C4864 raven_soc_0|gpio_outenb<1> BU_3VX2_71|Q 0.43fF
C4865 BU_3VX2_31|A raven_soc_0|gpio_out<8> 0.01fF
C4866 BU_3VX2_29|A raven_soc_0|flash_io3_di 3.46fF
C4867 IN_3VX2_1|A apllc03_1v8_0|B_CP 4.73fF
C4868 IN_3VX2_1|A LS_3VX2_15|A 0.01fF
C4869 raven_soc_0|gpio_out<7> vdd 0.34fF
C4870 VDD raven_padframe_0|FILLER20F_3|GNDO 0.07fF
C4871 AMUX2_3V_0|SEL BU_3VX2_54|Q 0.08fF
C4872 raven_soc_0|gpio_outenb<12> BU_3VX2_24|Q 0.01fF
C4873 raven_soc_0|gpio_pullup<15> BU_3VX2_27|Q 0.01fF
C4874 raven_soc_0|gpio_outenb<11> BU_3VX2_23|Q 0.01fF
C4875 raven_soc_0|gpio_outenb<15> BU_3VX2_26|Q 0.01fF
C4876 raven_soc_0|gpio_outenb<14> BU_3VX2_25|Q 0.01fF
C4877 raven_soc_0|gpio_outenb<6> apllc03_1v8_0|CLK 0.01fF
C4878 BU_3VX2_24|A BU_3VX2_63|A 0.01fF
C4879 BU_3VX2_10|A BU_3VX2_3|A 1.57fF
C4880 BU_3VX2_9|A BU_3VX2_4|A 2.47fF
C4881 BU_3VX2_10|A BU_3VX2_15|A 2.64fF
C4882 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<11> 0.12fF
C4883 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<7> 0.01fF
C4884 BU_3VX2_37|A raven_soc_0|flash_io3_di 0.01fF
C4885 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<4> 0.54fF
C4886 BU_3VX2_35|A raven_soc_0|flash_io1_oeb 0.01fF
C4887 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<9> 19.17fF
C4888 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<0> 0.01fF
C4889 AMUX4_3V_4|AOUT raven_soc_0|flash_clk 6.74fF
C4890 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<7> 0.01fF
C4891 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<9> 0.01fF
C4892 raven_soc_0|ext_clk raven_soc_0|flash_io3_do 34.56fF
C4893 raven_soc_0|gpio_in<7> raven_soc_0|gpio_in<11> 7.35fF
C4894 raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<15> 10.56fF
C4895 AMUX4_3V_3|SEL[1] AMUX4_3V_3|SEL[0] 189.35fF
C4896 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<10> 18.40fF
C4897 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_out<15> 0.02fF
C4898 raven_soc_0|ext_clk AMUX4_3V_4|AIN3 17.50fF
C4899 LS_3VX2_15|Q LS_3VX2_17|Q 4.68fF
C4900 BU_3VX2_61|A BU_3VX2_62|A 1.25fF
C4901 BU_3VX2_49|Q vdd 2.75fF
C4902 AMUX4_3V_0|SEL[0] BU_3VX2_50|Q 8.83fF
C4903 BU_3VX2_3|A BU_3VX2_0|A 0.01fF
C4904 BU_3VX2_0|A BU_3VX2_15|A 0.01fF
C4905 BU_3VX2_22|A BU_3VX2_31|A 2.37fF
C4906 raven_padframe_0|APR00DF_5|VDDO raven_padframe_0|APR00DF_5|GNDO 2.28fF
C4907 raven_padframe_0|FILLER20F_4|GNDR raven_padframe_0|FILLER20F_4|GNDO 0.81fF
C4908 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_in<3> 1.76fF
C4909 raven_spi_0|sdo_enb LOGIC0_3V_3|Q 2.05fF
C4910 BU_3VX2_65|A BU_3VX2_33|A 2.01fF
C4911 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<12> 0.22fF
C4912 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<7> 0.20fF
C4913 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<10> 0.61fF
C4914 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<7> 0.01fF
C4915 markings_0|efabless_logo_0|m1_7500_n8250# markings_0|efabless_logo_0|m1_6600_n9150# 0.33fF
C4916 markings_0|efabless_logo_0|m1_2700_n10050# markings_0|efabless_logo_0|m1_4500_n11550# 0.01fF
C4917 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<7> 3.25fF
C4918 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<25> 0.01fF
C4919 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<12> 3.88fF
C4920 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<14> 19.25fF
C4921 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<0> 0.11fF
C4922 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<15> 15.16fF
C4923 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<13> 16.74fF
C4924 raven_soc_0|gpio_out<14> raven_soc_0|ext_clk 0.01fF
C4925 raven_soc_0|gpio_in<5> raven_soc_0|gpio_pullup<5> 0.30fF
C4926 raven_soc_0|gpio_outenb<8> VDD3V3 0.07fF
C4927 LS_3VX2_19|A LS_3VX2_16|A 53.76fF
C4928 raven_soc_0|ram_rdata<5> vdd 0.80fF
C4929 BU_3VX2_58|Q BU_3VX2_57|Q 232.62fF
C4930 BU_3VX2_60|Q BU_3VX2_55|Q 27.92fF
C4931 LS_3VX2_16|A BU_3VX2_52|Q 7.84fF
C4932 BU_3VX2_59|Q BU_3VX2_56|Q 50.78fF
C4933 BU_3VX2_61|Q BU_3VX2_54|Q 18.45fF
C4934 raven_padframe_0|VDDPADF_0|VDDR raven_padframe_0|VDDPADF_0|GNDO 0.13fF
C4935 BU_3VX2_25|A BU_3VX2_14|A 1.82fF
C4936 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<0> 0.01fF
C4937 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<8> 1.40fF
C4938 LS_3VX2_22|Q VDD3V3 2.51fF
C4939 VDD raven_padframe_0|CORNERESDF_3|GNDR 0.16fF
C4940 IN_3VX2_1|Q BU_3VX2_42|Q 0.01fF
C4941 BU_3VX2_12|A raven_soc_0|flash_io2_do 0.01fF
C4942 LS_3VX2_4|Q vdd 0.01fF
C4943 BU_3VX2_0|Q BU_3VX2_38|Q 0.01fF
C4944 BU_3VX2_0|Q BU_3VX2_67|Q 0.01fF
C4945 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_outenb<13> 0.03fF
C4946 raven_soc_0|gpio_pulldown<3> BU_3VX2_71|Q 0.23fF
C4947 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<24> 0.08fF
C4948 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<7> 15.27fF
C4949 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<30> 0.88fF
C4950 raven_soc_0|ram_rdata<4> raven_soc_0|ram_addr<3> 0.04fF
C4951 raven_soc_0|ram_rdata<24> raven_soc_0|ram_addr<4> 4.48fF
C4952 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<6> 48.95fF
C4953 raven_soc_0|ram_rdata<18> raven_soc_0|ram_addr<2> 0.07fF
C4954 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<9> 2.84fF
C4955 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<20> 0.01fF
C4956 BU_3VX2_37|Q BU_3VX2_70|Q 0.01fF
C4957 BU_3VX2_47|Q BU_3VX2_72|Q 2.01fF
C4958 raven_padframe_0|axtoc02_3v3_0|VDDR raven_padframe_0|axtoc02_3v3_0|VDDO 0.09fF
C4959 markings_0|manufacturer_0|_alphabet_L_0|m2_0_0# markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# 1.08fF
C4960 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<6> 5.89fF
C4961 LS_3VX2_3|Q raven_soc_0|flash_io3_di 0.01fF
C4962 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<9> 0.45fF
C4963 IN_3VX2_1|A AMUX4_3V_1|SEL[1] 0.01fF
C4964 IN_3VX2_1|A raven_soc_0|flash_io1_do 5.21fF
C4965 adc_low LS_3VX2_16|A 0.05fF
C4966 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<6> 0.08fF
C4967 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<15> 1.03fF
C4968 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<11> 0.28fF
C4969 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<8> 1.07fF
C4970 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<12> 11.97fF
C4971 BU_3VX2_0|Q raven_soc_0|flash_io1_oeb 0.28fF
C4972 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<15> 0.02fF
C4973 acsoc01_3v3_0|CS2_200N acsoc01_3v3_0|CS3_200N 0.04fF
C4974 raven_soc_0|gpio_in<1> BU_3VX2_71|Q 0.34fF
C4975 BU_3VX2_63|A BU_3VX2_16|A 0.01fF
C4976 BU_3VX2_4|A BU_3VX2_28|A 0.01fF
C4977 BU_3VX2_7|A BU_3VX2_27|A 0.01fF
C4978 BU_3VX2_63|A BU_3VX2_29|A 0.01fF
C4979 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<1> 2.90fF
C4980 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<10> 0.20fF
C4981 BU_3VX2_31|A raven_soc_0|gpio_pulldown<2> 0.01fF
C4982 LOGIC0_3V_4|Q raven_soc_0|flash_io3_di 0.08fF
C4983 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<8> 3.22fF
C4984 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_outenb<13> 13.69fF
C4985 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<14> 0.03fF
C4986 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<8> 6.06fF
C4987 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<10> 8.39fF
C4988 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pullup<13> 29.91fF
C4989 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<5> 0.01fF
C4990 raven_soc_0|gpio_outenb<5> BU_3VX2_71|Q 0.01fF
C4991 raven_soc_0|gpio_out<7> raven_soc_0|gpio_outenb<9> 2.54fF
C4992 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<13> 0.02fF
C4993 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<26> 0.36fF
C4994 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<27> 0.80fF
C4995 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<29> 0.61fF
C4996 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<3> 5.17fF
C4997 BU_3VX2_6|Q BU_3VX2_15|Q 8.83fF
C4998 BU_3VX2_2|Q BU_3VX2_69|Q 0.01fF
C4999 BU_3VX2_66|Q BU_3VX2_65|Q 20.70fF
C5000 BU_3VX2_15|Q BU_3VX2_7|Q 4.49fF
C5001 BU_3VX2_16|Q BU_3VX2_38|Q 1.14fF
C5002 BU_3VX2_19|Q BU_3VX2_22|Q 13.11fF
C5003 BU_3VX2_21|Q BU_3VX2_31|Q 2.87fF
C5004 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<2> 1.04fF
C5005 BU_3VX2_16|Q BU_3VX2_67|Q 0.05fF
C5006 BU_3VX2_6|Q BU_3VX2_9|Q 15.15fF
C5007 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<21> 0.38fF
C5008 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<19> 5.79fF
C5009 BU_3VX2_18|Q BU_3VX2_22|Q 11.23fF
C5010 BU_3VX2_5|Q BU_3VX2_17|Q 2.69fF
C5011 BU_3VX2_7|Q BU_3VX2_9|Q 24.57fF
C5012 BU_3VX2_30|Q BU_3VX2_67|Q 0.58fF
C5013 BU_3VX2_65|Q BU_3VX2_20|Q 0.02fF
C5014 LS_3VX2_22|A BU_3VX2_57|Q 0.02fF
C5015 BU_3VX2_40|Q vdd 2.44fF
C5016 raven_padframe_0|POWERCUTVDD3FC_1|GNDR raven_padframe_0|POWERCUTVDD3FC_1|VDDO 0.09fF
C5017 BU_3VX2_37|A BU_3VX2_63|A 0.01fF
C5018 BU_3VX2_21|A BU_3VX2_31|A 2.08fF
C5019 LS_3VX2_14|A AMUX2_3V_0|SEL 163.96fF
C5020 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<8> 0.01fF
C5021 BU_3VX2_64|A BU_3VX2_69|A 2.47fF
C5022 raven_padframe_0|VDDORPADF_3|GNDR raven_padframe_0|VDDORPADF_3|GNDO 0.81fF
C5023 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<15> 16.08fF
C5024 BU_3VX2_63|Q raven_soc_0|gpio_outenb<0> 0.01fF
C5025 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<9> 1.00fF
C5026 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<7> 0.01fF
C5027 BU_3VX2_73|Q adc0_data<5> 7.87fF
C5028 AMUX4_3V_3|SEL[1] BU_3VX2_26|Q 0.21fF
C5029 raven_soc_0|ram_rdata<13> vdd 0.82fF
C5030 raven_soc_0|ram_wdata<25> apllc03_1v8_0|CLK 0.01fF
C5031 raven_soc_0|gpio_in<14> raven_padframe_0|BBCUD4F_14|PO 0.04fF
C5032 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_in<4> 0.31fF
C5033 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<9> 0.08fF
C5034 LS_3VX2_9|Q LS_3VX2_24|Q 0.01fF
C5035 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<12> 0.06fF
C5036 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<15> 0.01fF
C5037 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<13> 0.63fF
C5038 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<12> 1.31fF
C5039 VDD raven_soc_0|irq_pin 0.17fF
C5040 BU_3VX2_8|A raven_soc_0|ext_clk 0.01fF
C5041 BU_3VX2_40|A BU_3VX2_40|Q 0.08fF
C5042 raven_padframe_0|FILLER20F_8|VDDR raven_padframe_0|FILLER20F_8|GNDO 0.13fF
C5043 raven_soc_0|gpio_in<2> BU_3VX2_40|Q 0.01fF
C5044 raven_soc_0|gpio_pulldown<1> raven_soc_0|ext_clk 0.01fF
C5045 raven_spi_0|sdo_enb VDD3V3 0.19fF
C5046 VDD raven_padframe_0|FILLER02F_1|GNDO 0.07fF
C5047 raven_soc_0|flash_io0_oeb raven_soc_0|flash_clk 394.42fF
C5048 raven_soc_0|flash_io0_di raven_soc_0|flash_io0_do 27.71fF
C5049 raven_soc_0|flash_io3_di raven_soc_0|flash_io1_oeb 26.12fF
C5050 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<31> 0.70fF
C5051 raven_padframe_0|APR00DF_0|VDDR raven_padframe_0|APR00DF_0|VDDO 0.06fF
C5052 BU_3VX2_1|Q LS_3VX2_23|A 6.08fF
C5053 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<17> 4.55fF
C5054 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<13> 4.29fF
C5055 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<15> 0.05fF
C5056 raven_soc_0|flash_io1_di raven_soc_0|ram_rdata<11> 1.15fF
C5057 raven_soc_0|ram_wdata<20> raven_soc_0|ram_addr<0> 0.01fF
C5058 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<16> 4.06fF
C5059 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<1> 0.01fF
C5060 LS_3VX2_16|A BU_3VX2_58|Q 16.78fF
C5061 raven_padframe_0|FILLER20F_3|GNDR raven_padframe_0|FILLER20F_3|GNDO 0.81fF
C5062 AMUX4_3V_3|AOUT AMUX4_3V_4|AIN2 0.84fF
C5063 BU_3VX2_9|A raven_soc_0|flash_io0_oeb 0.01fF
C5064 BU_3VX2_19|A raven_soc_0|flash_io3_oeb 0.01fF
C5065 BU_3VX2_3|A vdd 0.23fF
C5066 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<3> 7.40fF
C5067 LOGIC0_3V_4|Q raven_soc_0|irq_pin 0.08fF
C5068 raven_padframe_0|ICF_2|VDDR raven_padframe_0|ICF_2|VDDO 0.06fF
C5069 LS_3VX2_14|A BU_3VX2_61|Q 0.01fF
C5070 BU_3VX2_31|A raven_soc_0|gpio_pulldown<6> 0.01fF
C5071 BU_3VX2_15|A vdd 0.06fF
C5072 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<14> 0.64fF
C5073 BU_3VX2_14|A BU_3VX2_13|Q 0.16fF
C5074 AMUX2_3V_0|SEL BU_3VX2_56|Q 0.12fF
C5075 raven_soc_0|gpio_outenb<7> vdd 0.29fF
C5076 raven_soc_0|gpio_pullup<9> BU_3VX2_28|Q 0.01fF
C5077 raven_soc_0|gpio_pullup<15> BU_3VX2_25|Q 0.01fF
C5078 raven_soc_0|gpio_pullup<11> BU_3VX2_23|Q 0.01fF
C5079 raven_soc_0|gpio_pullup<8> apllc03_1v8_0|CLK 0.01fF
C5080 raven_soc_0|gpio_pullup<12> BU_3VX2_24|Q 0.01fF
C5081 BU_3VX2_63|A LS_3VX2_3|Q 0.23fF
C5082 IN_3VX2_1|Q adc_high 0.26fF
C5083 BU_3VX2_18|A BU_3VX2_26|A 2.71fF
C5084 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<11> 0.01fF
C5085 raven_soc_0|gpio_pulldown<13> BU_3VX2_0|Q 0.01fF
C5086 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<9> 20.44fF
C5087 LS_3VX2_3|A raven_soc_0|gpio_pullup<3> 0.01fF
C5088 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<9> 0.01fF
C5089 BU_3VX2_25|A raven_soc_0|flash_io1_do 0.01fF
C5090 BU_3VX2_63|Q raven_soc_0|flash_io0_do 0.01fF
C5091 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<8> 1.39fF
C5092 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<13> 0.84fF
C5093 raven_soc_0|gpio_in<15> VDD3V3 2.98fF
C5094 BU_3VX2_40|Q raven_soc_0|gpio_in<11> 0.01fF
C5095 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<6> 1.94fF
C5096 BU_3VX2_53|A LS_3VX2_16|Q 0.12fF
C5097 BU_3VX2_56|A BU_3VX2_60|A 0.76fF
C5098 BU_3VX2_57|A BU_3VX2_59|A 2.55fF
C5099 BU_3VX2_54|A LS_3VX2_15|Q 0.17fF
C5100 BU_3VX2_55|A BU_3VX2_61|A 0.38fF
C5101 BU_3VX2_52|A LS_3VX2_17|Q 0.09fF
C5102 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<3> 2.69fF
C5103 AMUX4_3V_0|SEL[0] BU_3VX2_48|Q 11.26fF
C5104 VDD3V3 BU_3VX2_43|Q 1.46fF
C5105 BU_3VX2_3|A BU_3VX2_40|A 1.43fF
C5106 LS_3VX2_9|A LS_3VX2_14|Q 0.16fF
C5107 LS_3VX2_6|Q LS_3VX2_9|Q 1.62fF
C5108 LS_3VX2_10|Q LS_3VX2_5|Q 9.55fF
C5109 BU_3VX2_18|A BU_3VX2_11|A 2.51fF
C5110 BU_3VX2_4|A BU_3VX2_14|A 1.03fF
C5111 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<13> 10.45fF
C5112 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_in<0> 48.81fF
C5113 BU_3VX2_66|A BU_3VX2_69|A 4.86fF
C5114 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<5> 1.52fF
C5115 BU_3VX2_31|A raven_soc_0|gpio_outenb<11> 0.01fF
C5116 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<0> 8.18fF
C5117 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<4> 0.28fF
C5118 raven_soc_0|gpio_pullup<1> BU_3VX2_0|Q 0.05fF
C5119 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<7> 0.01fF
C5120 raven_soc_0|gpio_outenb<9> BU_3VX2_40|Q 0.22fF
C5121 raven_soc_0|gpio_out<10> raven_soc_0|gpio_pullup<5> 0.02fF
C5122 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<14> 44.70fF
C5123 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<8> 2.50fF
C5124 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<0> 0.04fF
C5125 raven_soc_0|flash_io1_oeb raven_soc_0|irq_pin 0.01fF
C5126 BU_3VX2_2|Q BU_3VX2_29|Q 0.96fF
C5127 BU_3VX2_21|Q apllc03_1v8_0|CLK 0.01fF
C5128 LS_3VX2_22|A LS_3VX2_16|A 0.01fF
C5129 BU_3VX2_10|Q BU_3VX2_29|Q 8.72fF
C5130 BU_3VX2_62|Q BU_3VX2_55|Q 18.45fF
C5131 BU_3VX2_22|Q BU_3VX2_27|Q 9.38fF
C5132 BU_3VX2_60|Q BU_3VX2_57|Q 49.46fF
C5133 BU_3VX2_17|Q BU_3VX2_28|Q 4.89fF
C5134 BU_3VX2_61|Q BU_3VX2_56|Q 27.14fF
C5135 LS_3VX2_15|A BU_3VX2_54|Q 12.04fF
C5136 BU_3VX2_8|Q apllc03_1v8_0|CLK 0.01fF
C5137 BU_3VX2_22|A BU_3VX2_21|A 39.08fF
C5138 LS_3VX2_8|Q LS_3VX2_9|Q 0.63fF
C5139 LS_3VX2_12|A LS_3VX2_8|A 152.41fF
C5140 BU_3VX2_23|A raven_soc_0|flash_csb 4.17fF
C5141 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<1> 11.65fF
C5142 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<14> 0.01fF
C5143 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<14> 0.01fF
C5144 raven_padframe_0|FILLER20FC_0|VDDR raven_padframe_0|FILLER20FC_0|VDDO 0.06fF
C5145 LS_3VX2_5|A BU_3VX2_55|Q 10.89fF
C5146 BU_3VX2_0|Q BU_3VX2_65|Q 0.01fF
C5147 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_pullup<13> 0.58fF
C5148 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_out<8> 3.26fF
C5149 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<14> 9.56fF
C5150 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<23> 0.03fF
C5151 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<8> 0.06fF
C5152 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<24> 0.41fF
C5153 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<4> 0.21fF
C5154 AMUX4_3V_3|SEL[1] BU_3VX2_11|Q 0.03fF
C5155 raven_soc_0|flash_io0_di raven_padframe_0|BBC4F_0|PO 0.04fF
C5156 raven_soc_0|flash_clk BU_3VX2_29|Q 12.42fF
C5157 raven_padframe_0|axtoc02_3v3_0|m4_0_22024# raven_padframe_0|axtoc02_3v3_0|VDDO 2.34fF
C5158 raven_soc_0|gpio_out<0> raven_soc_0|ext_clk 0.01fF
C5159 BU_3VX2_63|A raven_soc_0|flash_io1_oeb 0.01fF
C5160 VDD raven_padframe_0|BBCUD4F_15|GNDR 0.16fF
C5161 IN_3VX2_1|A raven_soc_0|gpio_in<10> 0.01fF
C5162 analog_out raven_soc_0|ser_tx 3.31fF
C5163 VDD raven_padframe_0|FILLER50F_1|GNDR 0.16fF
C5164 BU_3VX2_28|A raven_soc_0|flash_io0_oeb 8.09fF
C5165 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<6> 0.01fF
C5166 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<14> 0.03fF
C5167 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<7> 0.12fF
C5168 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<8> 0.21fF
C5169 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<11> 0.02fF
C5170 BU_3VX2_29|A BU_3VX2_26|Q 0.02fF
C5171 raven_soc_0|gpio_out<12> raven_soc_0|ext_clk 0.01fF
C5172 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pullup<5> 0.02fF
C5173 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<15> 9.60fF
C5174 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<5> 0.95fF
C5175 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<15> 0.02fF
C5176 raven_soc_0|gpio_out<13> VDD3V3 0.07fF
C5177 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<19> 4.39fF
C5178 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<23> 0.32fF
C5179 LOGIC1_3V_3|Q LOGIC1_3V_2|Q 0.58fF
C5180 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<14> 0.01fF
C5181 BU_3VX2_5|A raven_soc_0|flash_io0_do 0.01fF
C5182 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<10> 6.53fF
C5183 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<9> 5.55fF
C5184 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<8> 17.31fF
C5185 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pullup<14> 0.07fF
C5186 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pullup<13> 17.97fF
C5187 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<8> 0.02fF
C5188 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<14> 0.02fF
C5189 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pulldown<7> 0.02fF
C5190 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pullup<6> 0.03fF
C5191 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pulldown<6> 5.25fF
C5192 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<5> 0.01fF
C5193 raven_soc_0|gpio_pullup<7> BU_3VX2_71|Q 0.01fF
C5194 BU_3VX2_35|Q BU_3VX2_15|Q 0.02fF
C5195 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<25> 1.10fF
C5196 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<12> 2.19fF
C5197 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<2> 0.01fF
C5198 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<14> 0.36fF
C5199 BU_3VX2_12|Q BU_3VX2_68|Q 3.13fF
C5200 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<25> 0.22fF
C5201 BU_3VX2_6|Q BU_3VX2_64|Q 0.02fF
C5202 BU_3VX2_35|Q BU_3VX2_9|Q 2.45fF
C5203 BU_3VX2_19|Q BU_3VX2_31|Q 2.22fF
C5204 BU_3VX2_31|Q BU_3VX2_18|Q 2.05fF
C5205 BU_3VX2_65|Q BU_3VX2_30|Q 0.53fF
C5206 BU_3VX2_64|Q BU_3VX2_7|Q 0.01fF
C5207 BU_3VX2_69|Q BU_3VX2_33|Q 0.55fF
C5208 VDD3V3 BU_3VX2_50|Q 0.15fF
C5209 BU_3VX2_23|A BU_3VX2_20|A 7.88fF
C5210 raven_spi_0|SDO LOGIC0_3V_4|Q 0.80fF
C5211 IN_3VX2_1|Q IN_3VX2_1|A 185.21fF
C5212 LS_3VX2_12|A LS_3VX2_4|A 12.43fF
C5213 BU_3VX2_71|A BU_3VX2_26|A 0.01fF
C5214 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<8> 0.01fF
C5215 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<10> 0.01fF
C5216 raven_padframe_0|CORNERESDF_1|VDDR raven_padframe_0|CORNERESDF_1|GNDO 0.13fF
C5217 LOGIC0_3V_0|Q raven_spi_0|SDI 2.29fF
C5218 raven_soc_0|flash_io0_oeb BU_3VX2_33|Q 0.01fF
C5219 AMUX4_3V_1|SEL[1] BU_3VX2_54|Q 27.95fF
C5220 raven_soc_0|ram_addr<7> vdd 0.19fF
C5221 raven_soc_0|ram_rdata<26> apllc03_1v8_0|CLK 0.01fF
C5222 raven_soc_0|flash_io1_di raven_padframe_0|BBC4F_1|PO 0.04fF
C5223 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<10> 0.19fF
C5224 BU_3VX2_71|A BU_3VX2_11|A 0.01fF
C5225 IN_3VX2_1|A raven_soc_0|gpio_in<0> 0.01fF
C5226 LS_3VX2_6|A LS_3VX2_13|A 18.16fF
C5227 IN_3VX2_1|A raven_soc_0|flash_csb 64.58fF
C5228 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<11> 0.01fF
C5229 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<12> 0.01fF
C5230 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<14> 0.01fF
C5231 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<13> 0.29fF
C5232 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<5> 1.08fF
C5233 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<9> 0.02fF
C5234 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<12> 7.80fF
C5235 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<7> 0.01fF
C5236 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<6> 0.01fF
C5237 LS_3VX2_10|A VDD3V3 0.51fF
C5238 BU_3VX2_18|A VDD3V3 0.39fF
C5239 LS_3VX2_7|A BU_3VX2_54|Q 7.54fF
C5240 raven_soc_0|ser_rx raven_soc_0|irq_pin 110.92fF
C5241 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<31> 8.67fF
C5242 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<20> 0.01fF
C5243 raven_soc_0|flash_io1_di raven_soc_0|flash_io0_di 391.84fF
C5244 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<16> 15.67fF
C5245 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<17> 19.94fF
C5246 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<13> 5.09fF
C5247 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<21> 33.43fF
C5248 BU_3VX2_36|Q BU_3VX2_20|Q 0.01fF
C5249 raven_soc_0|ram_rdata<21> raven_soc_0|ram_addr<0> 4.70fF
C5250 BU_3VX2_66|Q BU_3VX2_36|Q 3.70fF
C5251 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<1> 1.66fF
C5252 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<29> 9.33fF
C5253 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<31> 0.01fF
C5254 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<22> 0.01fF
C5255 raven_soc_0|flash_io2_do raven_soc_0|flash_clk 21.30fF
C5256 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<27> 0.01fF
C5257 LS_3VX2_16|A BU_3VX2_60|Q 25.99fF
C5258 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<4> 0.01fF
C5259 raven_spi_0|SDO raven_soc_0|flash_io1_oeb 0.39fF
C5260 raven_soc_0|gpio_pullup<2> BU_3VX2_40|Q 0.02fF
C5261 BU_3VX2_9|A raven_soc_0|flash_io2_do 0.01fF
C5262 LS_3VX2_13|Q LS_3VX2_19|A 0.01fF
C5263 LS_3VX2_14|A LS_3VX2_15|A 0.02fF
C5264 BU_3VX2_4|A raven_soc_0|flash_io1_do 0.01fF
C5265 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<6> 0.49fF
C5266 BU_3VX2_28|A BU_3VX2_29|Q 0.03fF
C5267 VDD raven_padframe_0|aregc01_3v3_0|VDDR 0.54fF
C5268 raven_soc_0|gpio_pullup<9> vdd 0.22fF
C5269 raven_soc_0|gpio_pulldown<9> BU_3VX2_28|Q 0.01fF
C5270 raven_soc_0|gpio_outenb<0> BU_3VX2_24|Q 0.01fF
C5271 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<9> 1.27fF
C5272 LS_3VX2_3|A raven_soc_0|gpio_pulldown<5> 0.01fF
C5273 BU_3VX2_14|A raven_soc_0|flash_io0_oeb 0.01fF
C5274 BU_3VX2_63|Q raven_soc_0|flash_io1_di 13.88fF
C5275 raven_soc_0|ext_clk raven_soc_0|gpio_pullup<5> 3.38fF
C5276 raven_soc_0|gpio_in<14> VDD3V3 0.07fF
C5277 BU_3VX2_52|A BU_3VX2_54|A 4.42fF
C5278 VDD3V3 BU_3VX2_56|A 0.05fF
C5279 LS_3VX2_20|A BU_3VX2_42|Q 158.50fF
C5280 raven_spi_0|SDI BU_3VX2_40|A 1.87fF
C5281 LS_3VX2_13|Q adc_low 0.12fF
C5282 BU_3VX2_20|A IN_3VX2_1|A 2.10fF
C5283 BU_3VX2_1|A BU_3VX2_65|A 0.51fF
C5284 BU_3VX2_31|A raven_soc_0|gpio_pullup<11> 0.01fF
C5285 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<7> 1.24fF
C5286 LS_3VX2_6|A raven_soc_0|ser_rx 0.01fF
C5287 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<9> 0.01fF
C5288 BU_3VX2_35|A BU_3VX2_71|Q 0.02fF
C5289 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<10> 0.01fF
C5290 markings_0|product_name_0|_alphabet_A_0|m2_0_0# markings_0|product_name_0|_alphabet_R_0|m2_0_0# 0.95fF
C5291 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<20> 0.21fF
C5292 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<0> 0.01fF
C5293 raven_soc_0|gpio_pulldown<15> BU_3VX2_71|Q 0.01fF
C5294 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<12> 0.02fF
C5295 raven_soc_0|gpio_pullup<6> VDD3V3 0.07fF
C5296 BU_3VX2_12|Q BU_3VX2_24|Q 4.31fF
C5297 BU_3VX2_15|Q BU_3VX2_23|Q 4.48fF
C5298 BU_3VX2_38|Q BU_3VX2_26|Q 0.01fF
C5299 BU_3VX2_19|Q apllc03_1v8_0|CLK 0.01fF
C5300 BU_3VX2_62|Q BU_3VX2_57|Q 24.88fF
C5301 BU_3VX2_9|Q BU_3VX2_23|Q 10.31fF
C5302 BU_3VX2_17|Q vdd 2.08fF
C5303 BU_3VX2_22|Q BU_3VX2_25|Q 14.56fF
C5304 LS_3VX2_15|A BU_3VX2_56|Q 16.53fF
C5305 BU_3VX2_31|Q BU_3VX2_27|Q 8.18fF
C5306 BU_3VX2_67|Q BU_3VX2_26|Q 0.01fF
C5307 BU_3VX2_18|Q apllc03_1v8_0|CLK 0.01fF
C5308 raven_padframe_0|BT4FC_0|VDDR LOGIC0_3V_4|Q 0.01fF
C5309 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<15> 0.01fF
C5310 LS_3VX2_5|A BU_3VX2_57|Q 8.56fF
C5311 raven_soc_0|ram_rdata<17> raven_soc_0|ram_addr<0> 0.72fF
C5312 raven_soc_0|ram_rdata<11> vdd 0.59fF
C5313 raven_soc_0|flash_io1_oeb BU_3VX2_26|Q 0.01fF
C5314 raven_soc_0|flash_io0_di BU_3VX2_28|Q 0.01fF
C5315 raven_soc_0|flash_io0_do BU_3VX2_24|Q 0.01fF
C5316 raven_soc_0|flash_io3_oeb BU_3VX2_27|Q 0.01fF
C5317 BU_3VX2_49|A vdd 0.06fF
C5318 raven_padframe_0|FILLER01F_1|GNDR raven_padframe_0|FILLER01F_1|GNDO 0.81fF
C5319 raven_padframe_0|FILLER50F_0|VDDR raven_padframe_0|FILLER50F_0|VDDO 0.06fF
C5320 raven_padframe_0|aregc01_3v3_1|VDDR raven_padframe_0|aregc01_3v3_1|VDDO 0.04fF
C5321 BU_3VX2_25|A raven_soc_0|flash_csb 4.78fF
C5322 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<9> 0.28fF
C5323 BU_3VX2_10|A raven_soc_0|flash_io0_di 0.06fF
C5324 BU_3VX2_5|A BU_3VX2_5|Q 0.08fF
C5325 LS_3VX2_14|A AMUX4_3V_1|SEL[1] 8.12fF
C5326 BU_3VX2_71|A VDD3V3 0.14fF
C5327 VDD raven_padframe_0|FILLER20F_8|GNDO 0.07fF
C5328 BU_3VX2_13|A BU_3VX2_12|Q 0.16fF
C5329 AMUX4_3V_4|AIN1 raven_soc_0|ser_tx 3.87fF
C5330 IN_3VX2_1|A raven_soc_0|gpio_in<13> 0.01fF
C5331 BU_3VX2_28|A raven_soc_0|flash_io2_do 3.74fF
C5332 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_in<9> 0.06fF
C5333 raven_soc_0|gpio_outenb<14> BU_3VX2_40|Q 0.32fF
C5334 LS_3VX2_3|A raven_soc_0|flash_io0_oeb 0.01fF
C5335 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<14> 0.02fF
C5336 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<15> 0.02fF
C5337 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<7> 0.01fF
C5338 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pullup<5> 0.02fF
C5339 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<6> 0.01fF
C5340 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<11> 7.92fF
C5341 raven_soc_0|gpio_outenb<12> raven_soc_0|ext_clk 0.01fF
C5342 raven_soc_0|gpio_outenb<15> VDD3V3 3.22fF
C5343 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<23> 0.10fF
C5344 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<19> 0.06fF
C5345 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<11> 6.28fF
C5346 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<20> 0.06fF
C5347 acmpc01_3v3_0|IBN BU_3VX2_32|A 12.68fF
C5348 LS_3VX2_14|A LS_3VX2_7|A 23.37fF
C5349 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<1> 45.67fF
C5350 LS_3VX2_12|A vdd 2.65fF
C5351 VDD raven_padframe_0|ICF_2|GNDO 0.07fF
C5352 BU_3VX2_5|A raven_soc_0|flash_io1_di 0.04fF
C5353 BU_3VX2_0|A raven_soc_0|flash_io0_di 28.07fF
C5354 BU_3VX2_13|A raven_soc_0|flash_io0_do 0.01fF
C5355 VDD raven_padframe_0|GNDORPADF_6|VDDR 0.71fF
C5356 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pullup<6> 8.71fF
C5357 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<9> 22.59fF
C5358 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<8> 0.02fF
C5359 BU_3VX2_33|A raven_soc_0|flash_io2_di 0.24fF
C5360 raven_soc_0|ram_wenb raven_soc_0|ram_addr<1> 0.01fF
C5361 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<2> 0.01fF
C5362 BU_3VX2_0|Q BU_3VX2_71|Q 105.30fF
C5363 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<14> 0.02fF
C5364 BU_3VX2_0|Q BU_3VX2_36|Q 0.01fF
C5365 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pulldown<6> 0.02fF
C5366 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<10> 0.01fF
C5367 raven_soc_0|gpio_pulldown<14> BU_3VX2_24|Q 0.01fF
C5368 BU_3VX2_63|Q BU_3VX2_28|Q 2.54fF
C5369 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<12> 0.01fF
C5370 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<2> 10.93fF
C5371 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<16> 2.74fF
C5372 raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<2> 14.51fF
C5373 BU_3VX2_68|Q BU_3VX2_5|Q 0.97fF
C5374 VDD3V3 LS_3VX2_27|Q 0.19fF
C5375 BU_3VX2_24|A BU_3VX2_26|A 19.42fF
C5376 VDD3V3 BU_3VX2_48|Q 0.02fF
C5377 raven_padframe_0|CORNERESDF_2|VDDR raven_padframe_0|CORNERESDF_2|VDDO 0.06fF
C5378 LS_3VX2_12|Q LS_3VX2_10|Q 1.59fF
C5379 raven_padframe_0|APR00DF_3|GNDR raven_padframe_0|APR00DF_3|VDDO 0.09fF
C5380 raven_padframe_0|FILLER02F_0|GNDR raven_padframe_0|FILLER02F_0|VDDO 0.09fF
C5381 raven_padframe_0|FILLER02F_1|GNDR raven_padframe_0|FILLER02F_1|GNDO 0.84fF
C5382 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<12> 0.01fF
C5383 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<13> 0.01fF
C5384 raven_soc_0|gpio_pulldown<0> BU_3VX2_71|Q 0.01fF
C5385 LOGIC0_3V_4|Q raven_padframe_0|ICFC_1|PO 0.04fF
C5386 BU_3VX2_1|Q raven_soc_0|ext_clk 2.23fF
C5387 raven_soc_0|ser_tx VDD3V3 3.50fF
C5388 raven_soc_0|ram_rdata<2> vdd 0.92fF
C5389 AMUX4_3V_1|SEL[1] BU_3VX2_56|Q 16.89fF
C5390 BU_3VX2_24|A BU_3VX2_11|A 1.60fF
C5391 BU_3VX2_53|A BU_3VX2_52|Q 0.03fF
C5392 raven_soc_0|irq_pin BU_3VX2_72|Q 0.02fF
C5393 VDD raven_padframe_0|BBCUD4F_9|VDDR 0.71fF
C5394 BU_3VX2_20|A BU_3VX2_25|A 4.41fF
C5395 LS_3VX2_9|Q LS_3VX2_14|Q 1.70fF
C5396 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<10> 0.01fF
C5397 BU_3VX2_31|A raven_soc_0|gpio_pulldown<8> 0.01fF
C5398 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<15> 0.01fF
C5399 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<3> 0.01fF
C5400 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<7> 0.01fF
C5401 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<6> 0.01fF
C5402 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<9> 0.15fF
C5403 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<14> 0.81fF
C5404 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<12> 10.80fF
C5405 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<15> 1.04fF
C5406 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<13> 0.02fF
C5407 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<12> 0.01fF
C5408 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<12> 13.48fF
C5409 LS_3VX2_19|Q VDD3V3 0.20fF
C5410 LS_3VX2_24|A VDD3V3 0.83fF
C5411 LS_3VX2_7|A BU_3VX2_56|Q 8.08fF
C5412 raven_padframe_0|BBCUD4F_7|VDDR raven_padframe_0|BBCUD4F_7|GNDR 0.68fF
C5413 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<9> 0.13fF
C5414 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<4> 22.73fF
C5415 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<31> 0.14fF
C5416 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<24> 1.94fF
C5417 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<20> 0.10fF
C5418 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<30> 7.20fF
C5419 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<21> 0.01fF
C5420 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<24> 0.01fF
C5421 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<23> 0.01fF
C5422 BU_3VX2_16|Q BU_3VX2_36|Q 0.41fF
C5423 raven_soc_0|flash_io3_do raven_soc_0|flash_io2_di 120.91fF
C5424 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io3_oeb 326.75fF
C5425 BU_3VX2_2|Q BU_3VX2_32|Q 0.01fF
C5426 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<13> 6.86fF
C5427 BU_3VX2_32|Q BU_3VX2_10|Q 1.39fF
C5428 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<2> 5.39fF
C5429 BU_3VX2_4|Q BU_3VX2_9|Q 11.71fF
C5430 BU_3VX2_70|Q BU_3VX2_17|Q 0.01fF
C5431 BU_3VX2_11|Q BU_3VX2_67|Q 0.61fF
C5432 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<15> 0.02fF
C5433 BU_3VX2_15|Q BU_3VX2_4|Q 4.59fF
C5434 BU_3VX2_36|Q BU_3VX2_30|Q 0.24fF
C5435 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<31> 4.00fF
C5436 BU_3VX2_38|Q BU_3VX2_11|Q 2.75fF
C5437 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<27> 2.87fF
C5438 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<22> 0.02fF
C5439 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<25> 2.23fF
C5440 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<26> 0.01fF
C5441 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<29> 0.01fF
C5442 raven_soc_0|flash_io1_do raven_soc_0|flash_io0_oeb 47.93fF
C5443 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<17> 0.01fF
C5444 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<21> 0.01fF
C5445 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<14> 5.40fF
C5446 LS_3VX2_16|A BU_3VX2_62|Q 169.51fF
C5447 BU_3VX2_45|A BU_3VX2_42|Q 0.02fF
C5448 AMUX4_3V_4|AIN2 BU_3VX2_59|Q 0.01fF
C5449 BU_3VX2_44|Q BU_3VX2_46|Q 83.21fF
C5450 BU_3VX2_42|Q BU_3VX2_47|Q 20.78fF
C5451 BU_3VX2_43|Q adc0_data<5> 32.87fF
C5452 BU_3VX2_29|Q apllc03_1v8_0|B_CP 4.17fF
C5453 apllc03_1v8_0|CLK BU_3VX2_27|Q 6.18fF
C5454 raven_padframe_0|BBCUD4F_9|VDDR LOGIC0_3V_4|Q 0.01fF
C5455 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<3> 1.34fF
C5456 BU_3VX2_2|A raven_soc_0|flash_io2_oeb 0.01fF
C5457 BU_3VX2_6|A raven_soc_0|flash_io3_oeb 0.01fF
C5458 LS_3VX2_13|Q LS_3VX2_22|A 0.01fF
C5459 LS_3VX2_11|A BU_3VX2_55|Q 7.58fF
C5460 IN_3VX2_1|Q BU_3VX2_54|Q 0.01fF
C5461 raven_padframe_0|FILLER50F_2|VDDR raven_padframe_0|FILLER50F_2|VDDO 0.06fF
C5462 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<3> 0.29fF
C5463 LS_3VX2_5|A LS_3VX2_16|A 0.01fF
C5464 raven_soc_0|gpio_pulldown<9> vdd 0.19fF
C5465 LS_3VX2_3|A BU_3VX2_29|Q 0.01fF
C5466 raven_soc_0|gpio_pulldown<10> BU_3VX2_24|Q 0.01fF
C5467 raven_soc_0|gpio_pulldown<13> BU_3VX2_26|Q 0.01fF
C5468 BU_3VX2_71|Q raven_soc_0|flash_io3_di 0.02fF
C5469 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<16> 11.97fF
C5470 raven_soc_0|flash_io1_oeb BU_3VX2_11|Q 0.06fF
C5471 BU_3VX2_6|A BU_3VX2_2|A 2.31fF
C5472 BU_3VX2_32|A BU_3VX2_70|A 0.55fF
C5473 BU_3VX2_65|A BU_3VX2_1|Q 0.02fF
C5474 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<7> 2.52fF
C5475 BU_3VX2_14|A raven_soc_0|flash_io2_do 0.01fF
C5476 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<15> 81.98fF
C5477 raven_soc_0|gpio_out<2> BU_3VX2_28|Q 0.01fF
C5478 raven_soc_0|gpio_outenb<2> BU_3VX2_23|Q 0.01fF
C5479 raven_soc_0|gpio_pullup<1> BU_3VX2_26|Q 0.01fF
C5480 BU_3VX2_44|A LS_3VX2_20|Q 0.81fF
C5481 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<0> 26.30fF
C5482 BU_3VX2_3|A BU_3VX2_7|A 3.10fF
C5483 BU_3VX2_10|A BU_3VX2_5|A 2.75fF
C5484 VDD raven_padframe_0|BBCUD4F_8|VDDR 0.71fF
C5485 raven_padframe_0|BT4F_1|GNDR raven_padframe_0|BT4F_1|GNDO 0.81fF
C5486 BU_3VX2_7|A BU_3VX2_15|A 1.44fF
C5487 BU_3VX2_17|A BU_3VX2_12|A 3.85fF
C5488 BU_3VX2_16|A BU_3VX2_26|A 2.09fF
C5489 IN_3VX2_1|A raven_soc_0|gpio_outenb<1> 0.01fF
C5490 BU_3VX2_29|A BU_3VX2_26|A 12.04fF
C5491 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<4> 1.11fF
C5492 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<2> 1.16fF
C5493 raven_soc_0|gpio_outenb<3> BU_3VX2_0|Q 0.01fF
C5494 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<9> 0.01fF
C5495 raven_padframe_0|BBCUD4F_1|GNDR raven_padframe_0|BBCUD4F_1|GNDO 0.81fF
C5496 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<12> 0.01fF
C5497 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<14> 37.83fF
C5498 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<8> 15.68fF
C5499 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<5> 0.01fF
C5500 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<14> 7.57fF
C5501 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_14|PO 0.04fF
C5502 raven_padframe_0|FILLER10F_0|VDDR raven_padframe_0|FILLER10F_0|GNDR 0.68fF
C5503 AMUX4_3V_3|SEL[1] VDD3V3 0.65fF
C5504 raven_soc_0|irq_pin AMUX4_3V_1|SEL[0] 0.01fF
C5505 BU_3VX2_31|Q BU_3VX2_25|Q 11.41fF
C5506 BU_3VX2_5|Q BU_3VX2_24|Q 1.39fF
C5507 BU_3VX2_68|Q BU_3VX2_28|Q 1.08fF
C5508 BU_3VX2_65|Q BU_3VX2_26|Q 1.13fF
C5509 BU_3VX2_64|Q BU_3VX2_23|Q 1.54fF
C5510 AMUX4_3V_4|SEL[1] apllc03_1v8_0|CLK 13.85fF
C5511 VDD raven_padframe_0|FILLER20F_5|VDDR 0.71fF
C5512 BU_3VX2_0|A BU_3VX2_5|A 0.05fF
C5513 raven_padframe_0|BBCUD4F_8|VDDR LOGIC0_3V_4|Q 0.01fF
C5514 BU_3VX2_37|A BU_3VX2_26|A 0.38fF
C5515 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<9> 0.28fF
C5516 BU_3VX2_16|A BU_3VX2_11|A 3.76fF
C5517 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<0> 2.68fF
C5518 BU_3VX2_4|A raven_soc_0|flash_csb 0.01fF
C5519 BU_3VX2_29|A BU_3VX2_11|A 0.01fF
C5520 raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<0> 7.96fF
C5521 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<17> 0.01fF
C5522 raven_soc_0|ram_wdata<25> raven_soc_0|ram_rdata<15> 1.07fF
C5523 raven_soc_0|ram_wdata<29> raven_soc_0|ram_rdata<17> 0.41fF
C5524 raven_soc_0|ram_wdata<31> raven_soc_0|ram_rdata<1> 15.79fF
C5525 raven_soc_0|ram_wdata<27> raven_soc_0|ram_rdata<13> 0.41fF
C5526 raven_soc_0|ram_wdata<21> raven_soc_0|ram_rdata<16> 0.07fF
C5527 raven_soc_0|ram_wdata<22> raven_soc_0|ram_addr<0> 0.01fF
C5528 raven_soc_0|flash_io0_di vdd 3.06fF
C5529 BU_3VX2_45|A BU_3VX2_42|A 0.28fF
C5530 raven_soc_0|flash_io3_oeb BU_3VX2_25|Q 0.01fF
C5531 BU_3VX2_58|A BU_3VX2_59|Q 0.15fF
C5532 raven_soc_0|flash_io1_di BU_3VX2_24|Q 0.01fF
C5533 raven_soc_0|flash_io2_oeb apllc03_1v8_0|CLK 0.01fF
C5534 LS_3VX2_16|Q BU_3VX2_60|Q 0.03fF
C5535 raven_soc_0|flash_io1_do BU_3VX2_29|Q 0.01fF
C5536 adc0_data<5> BU_3VX2_50|Q 39.62fF
C5537 BU_3VX2_46|Q vdd 1.79fF
C5538 BU_3VX2_37|A BU_3VX2_11|A 1.99fF
C5539 BU_3VX2_37|A LOGIC0_3V_3|Q 0.43fF
C5540 raven_padframe_0|FILLER20F_5|VDDR LOGIC0_3V_4|Q 0.01fF
C5541 raven_padframe_0|BBCUD4F_9|GNDR raven_padframe_0|BBCUD4F_9|VDDO 0.09fF
C5542 AMUX4_3V_4|AOUT raven_soc_0|flash_csb 6.43fF
C5543 raven_padframe_0|aregc01_3v3_1|m4_0_22024# raven_padframe_0|aregc01_3v3_1|VDDO 1.17fF
C5544 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<7> 0.61fF
C5545 raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# raven_padframe_0|axtoc02_3v3_0|m4_55000_28769# 0.22fF
C5546 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<6> 1.08fF
C5547 BU_3VX2_24|A VDD3V3 0.71fF
C5548 BU_3VX2_8|A BU_3VX2_7|Q 0.16fF
C5549 BU_3VX2_8|A BU_3VX2_6|Q 0.03fF
C5550 VDD raven_padframe_0|APR00DF_5|GNDR 0.16fF
C5551 IN_3VX2_1|A LS_3VX2_20|A 0.01fF
C5552 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<14> 0.02fF
C5553 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<11> 6.94fF
C5554 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<5> 0.50fF
C5555 raven_soc_0|gpio_pullup<15> BU_3VX2_40|Q 0.06fF
C5556 LS_3VX2_3|A raven_soc_0|flash_io2_do 0.01fF
C5557 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<9> 4.31fF
C5558 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<15> 0.02fF
C5559 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<10> 0.02fF
C5560 raven_soc_0|gpio_pullup<12> raven_soc_0|ext_clk 0.01fF
C5561 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<0> 3.62fF
C5562 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<23> 147.15fF
C5563 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<20> 52.42fF
C5564 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<11> 3.05fF
C5565 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<28> 0.03fF
C5566 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<19> 0.29fF
C5567 raven_soc_0|gpio_outenb<8> BU_3VX2_27|Q 0.01fF
C5568 BU_3VX2_8|A raven_soc_0|flash_io2_di 0.01fF
C5569 BU_3VX2_63|A BU_3VX2_71|Q 0.16fF
C5570 BU_3VX2_40|A raven_soc_0|flash_io0_di 0.86fF
C5571 LOGIC0_3V_4|Q raven_soc_0|gpio_in<8> 0.08fF
C5572 adc_low LS_3VX2_19|A 5.24fF
C5573 BU_3VX2_13|A raven_soc_0|flash_io1_di 0.01fF
C5574 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<6> 5.73fF
C5575 LS_3VX2_6|A AMUX4_3V_1|SEL[0] 15.15fF
C5576 raven_soc_0|gpio_in<2> raven_soc_0|flash_io0_di 0.33fF
C5577 BU_3VX2_0|Q raven_soc_0|gpio_pullup<14> 0.23fF
C5578 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<13> 70.74fF
C5579 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pulldown<6> 0.02fF
C5580 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<9> 36.61fF
C5581 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<16> 2.36fF
C5582 adc_low BU_3VX2_52|Q 0.05fF
C5583 BU_3VX2_27|A raven_soc_0|flash_io3_oeb 4.53fF
C5584 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<5> 0.01fF
C5585 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<2> 19.02fF
C5586 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<8> 6.25fF
C5587 AMUX2_3V_0|SEL AMUX4_3V_4|AIN2 6.18fF
C5588 BU_3VX2_63|Q vdd 0.18fF
C5589 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_5|PO 0.04fF
C5590 raven_padframe_0|FILLER20F_3|VDDR raven_padframe_0|FILLER20F_3|VDDO 0.06fF
C5591 BU_3VX2_20|A BU_3VX2_4|A 0.48fF
C5592 BU_3VX2_19|A BU_3VX2_18|A 36.68fF
C5593 BU_3VX2_2|A BU_3VX2_27|A 0.01fF
C5594 LS_3VX2_3|Q BU_3VX2_26|A 0.01fF
C5595 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<13> 0.01fF
C5596 raven_soc_0|ram_wdata<16> vdd 0.61fF
C5597 raven_soc_0|irq_pin LS_3VX2_17|A 0.01fF
C5598 raven_soc_0|ram_wdata<2> vdd 2.10fF
C5599 raven_soc_0|gpio_in<1> IN_3VX2_1|A 0.01fF
C5600 BU_3VX2_52|A BU_3VX2_53|Q 0.15fF
C5601 LS_3VX2_7|Q LS_3VX2_9|Q 0.91fF
C5602 LS_3VX2_11|Q LS_3VX2_5|Q 1.93fF
C5603 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<4> 0.01fF
C5604 LS_3VX2_3|Q BU_3VX2_11|A 0.01fF
C5605 BU_3VX2_40|A BU_3VX2_63|Q 0.16fF
C5606 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<11> 0.29fF
C5607 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<8> 0.33fF
C5608 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<5> 0.08fF
C5609 raven_soc_0|gpio_in<2> BU_3VX2_63|Q 0.01fF
C5610 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<15> 0.02fF
C5611 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<7> 0.05fF
C5612 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_out<9> 0.39fF
C5613 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<10> 5.60fF
C5614 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<11> 32.64fF
C5615 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<14> 0.02fF
C5616 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<12> 11.91fF
C5617 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<26> 2.71fF
C5618 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<2> 0.39fF
C5619 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<13> 0.02fF
C5620 raven_soc_0|flash_io2_do raven_soc_0|flash_io1_do 349.21fF
C5621 BU_3VX2_13|Q BU_3VX2_14|Q 69.71fF
C5622 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<1> 0.06fF
C5623 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<4> 0.38fF
C5624 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<5> 0.46fF
C5625 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<7> 8.47fF
C5626 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<14> 4.11fF
C5627 BU_3VX2_15|Q BU_3VX2_3|Q 4.21fF
C5628 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<2> 0.58fF
C5629 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<17> 1.39fF
C5630 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<30> 0.76fF
C5631 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<21> 0.04fF
C5632 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<10> 0.06fF
C5633 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<8> 12.30fF
C5634 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<12> 0.31fF
C5635 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<21> 10.19fF
C5636 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<6> 0.11fF
C5637 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<19> 0.23fF
C5638 raven_soc_0|gpio_out<15> raven_soc_0|flash_io1_di 0.65fF
C5639 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<14> 0.01fF
C5640 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<24> 3.40fF
C5641 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<2> 0.01fF
C5642 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<4> 0.01fF
C5643 BU_3VX2_4|Q BU_3VX2_64|Q 2.70fF
C5644 BU_3VX2_3|Q BU_3VX2_9|Q 6.33fF
C5645 BU_3VX2_32|Q BU_3VX2_33|Q 0.57fF
C5646 AMUX4_3V_4|AIN2 BU_3VX2_61|Q 0.01fF
C5647 BU_3VX2_24|Q BU_3VX2_28|Q 69.86fF
C5648 BU_3VX2_23|Q apllc03_1v8_0|B_VCO 0.81fF
C5649 BU_3VX2_25|Q apllc03_1v8_0|CLK 1.40fF
C5650 LOGIC0_3V_4|Q LOGIC0_3V_3|Q 0.43fF
C5651 raven_padframe_0|CORNERESDF_0|GNDR raven_padframe_0|CORNERESDF_0|VDDO 0.09fF
C5652 LOGIC0_3V_4|Q raven_soc_0|gpio_out<5> 0.01fF
C5653 raven_soc_0|gpio_out<1> LS_3VX2_3|A 0.01fF
C5654 IN_3VX2_1|Q BU_3VX2_56|Q 0.01fF
C5655 BU_3VX2_38|A raven_soc_0|flash_io3_do 0.01fF
C5656 BU_3VX2_16|A VDD3V3 0.48fF
C5657 raven_padframe_0|FILLER20F_1|VDDR raven_padframe_0|FILLER20F_1|GNDR 0.68fF
C5658 LS_3VX2_11|A BU_3VX2_57|Q 6.34fF
C5659 BU_3VX2_29|A VDD3V3 1.37fF
C5660 raven_soc_0|gpio_pulldown<12> BU_3VX2_24|Q 0.01fF
C5661 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<13> 1.27fF
C5662 LS_3VX2_19|A BU_3VX2_58|Q 10.91fF
C5663 BU_3VX2_58|Q BU_3VX2_52|Q 22.11fF
C5664 BU_3VX2_37|A VDD3V3 0.32fF
C5665 VDD raven_padframe_0|FILLER01F_1|GNDO 0.07fF
C5666 BU_3VX2_5|A vdd 0.14fF
C5667 BU_3VX2_26|A raven_soc_0|flash_io1_oeb 3.59fF
C5668 raven_soc_0|gpio_out<3> BU_3VX2_40|Q 0.01fF
C5669 LS_3VX2_6|A LS_3VX2_17|A 0.09fF
C5670 BU_3VX2_63|Q raven_soc_0|gpio_in<11> 0.28fF
C5671 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<9> 0.01fF
C5672 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<6> 0.01fF
C5673 BU_3VX2_0|Q raven_soc_0|ram_wdata<23> 0.02fF
C5674 raven_soc_0|gpio_out<2> vdd 0.19fF
C5675 BU_3VX2_10|A BU_3VX2_13|A 4.71fF
C5676 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<7> 0.01fF
C5677 analog_out raven_soc_0|ser_rx 3.78fF
C5678 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<3> 0.97fF
C5679 AMUX4_3V_3|AOUT raven_soc_0|flash_clk 9.16fF
C5680 BU_3VX2_11|A raven_soc_0|flash_io1_oeb 0.01fF
C5681 raven_soc_0|gpio_in<3> raven_soc_0|flash_io0_do 7.10fF
C5682 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<6> 4.84fF
C5683 BU_3VX2_63|Q raven_soc_0|gpio_outenb<9> 0.33fF
C5684 IN_3VX2_1|A BU_3VX2_47|Q 6.80fF
C5685 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<10> 0.01fF
C5686 adc_low BU_3VX2_58|Q 0.05fF
C5687 raven_soc_0|flash_csb raven_soc_0|flash_io0_oeb 145.04fF
C5688 BU_3VX2_73|Q AMUX4_3V_0|SEL[1] 0.32fF
C5689 BU_3VX2_68|Q vdd 0.70fF
C5690 BU_3VX2_73|Q BU_3VX2_51|Q 14.95fF
C5691 raven_padframe_0|FILLER20FC_0|VDDR LOGIC0_3V_4|Q 0.01fF
C5692 BU_3VX2_19|A BU_3VX2_71|A 0.01fF
C5693 BU_3VX2_5|A BU_3VX2_40|A 0.93fF
C5694 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<9> 0.01fF
C5695 BU_3VX2_0|A BU_3VX2_13|A 0.01fF
C5696 BU_3VX2_31|A raven_soc_0|gpio_outenb<2> 0.01fF
C5697 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<2> 39.60fF
C5698 raven_soc_0|ram_addr<8> raven_soc_0|ram_addr<9> 63.04fF
C5699 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<13> 0.05fF
C5700 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<15> 4.87fF
C5701 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<0> 11.11fF
C5702 LS_3VX2_22|A LS_3VX2_19|A 41.86fF
C5703 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<17> 5.66fF
C5704 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<29> 0.01fF
C5705 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<31> 0.01fF
C5706 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<22> 0.01fF
C5707 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<27> 0.01fF
C5708 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<16> 1.41fF
C5709 raven_soc_0|ram_wdata<22> raven_soc_0|ram_wdata<29> 15.48fF
C5710 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<15> 0.64fF
C5711 LS_3VX2_22|A BU_3VX2_52|Q 0.02fF
C5712 raven_soc_0|ram_wdata<19> raven_soc_0|ram_rdata<1> 0.07fF
C5713 raven_soc_0|ram_wdata<26> raven_soc_0|ram_rdata<13> 0.02fF
C5714 BU_3VX2_47|A BU_3VX2_44|A 0.76fF
C5715 BU_3VX2_49|A LS_3VX2_21|Q 0.13fF
C5716 BU_3VX2_48|A LS_3VX2_20|Q 0.19fF
C5717 BU_3VX2_50|A BU_3VX2_42|A 0.13fF
C5718 LS_3VX2_16|Q BU_3VX2_62|Q 1.07fF
C5719 raven_soc_0|gpio_out<15> BU_3VX2_28|Q 0.01fF
C5720 raven_soc_0|gpio_in<10> BU_3VX2_29|Q 0.01fF
C5721 raven_soc_0|flash_io3_do BU_3VX2_23|Q 0.01fF
C5722 raven_soc_0|gpio_in<15> BU_3VX2_27|Q 0.01fF
C5723 BU_3VX2_58|A BU_3VX2_61|Q 0.02fF
C5724 adc0_data<5> BU_3VX2_48|Q 78.18fF
C5725 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<11> 0.01fF
C5726 raven_padframe_0|aregc01_3v3_1|m4_92500_30653# raven_padframe_0|aregc01_3v3_1|VDDR 0.07fF
C5727 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<7> 0.01fF
C5728 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<14> 0.01fF
C5729 raven_padframe_0|axtoc02_3v3_0|m4_55000_30653# raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# 0.17fF
C5730 raven_padframe_0|axtoc02_3v3_0|m4_0_29057# raven_padframe_0|axtoc02_3v3_0|m4_0_22024# 0.03fF
C5731 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<11> 4.05fF
C5732 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<12> 56.40fF
C5733 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<9> 0.01fF
C5734 VDD VDD3V3 4.00fF
C5735 BU_3VX2_18|A BU_3VX2_19|Q 0.03fF
C5736 BU_3VX2_18|A BU_3VX2_18|Q 0.08fF
C5737 LS_3VX2_3|Q VDD3V3 0.77fF
C5738 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<8> 0.01fF
C5739 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<5> 0.22fF
C5740 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<13> 0.02fF
C5741 BU_3VX2_0|Q raven_soc_0|gpio_in<9> 0.01fF
C5742 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<15> 8.72fF
C5743 raven_soc_0|gpio_outenb<0> raven_soc_0|ext_clk 0.01fF
C5744 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<6> 0.01fF
C5745 raven_soc_0|gpio_out<14> BU_3VX2_23|Q 0.01fF
C5746 BU_3VX2_71|Q BU_3VX2_26|Q 2.21fF
C5747 BU_3VX2_36|Q BU_3VX2_26|Q 0.01fF
C5748 BU_3VX2_23|A BU_3VX2_20|Q 0.02fF
C5749 BU_3VX2_20|A raven_soc_0|flash_io0_oeb 0.01fF
C5750 VDD raven_padframe_0|VDDORPADF_4|GNDR 0.16fF
C5751 LS_3VX2_11|A LS_3VX2_16|A 0.01fF
C5752 raven_spi_0|sdo_enb raven_soc_0|flash_io2_oeb 0.52fF
C5753 LOGIC0_3V_4|Q VDD3V3 9.34fF
C5754 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<13> 217.74fF
C5755 adc_low LS_3VX2_22|A 7.71fF
C5756 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pulldown<3> 20.57fF
C5757 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<11> 0.09fF
C5758 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pulldown<7> 0.02fF
C5759 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<5> 0.01fF
C5760 LS_3VX2_24|A adc0_data<5> 5.19fF
C5761 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<10> 26.07fF
C5762 raven_padframe_0|FILLER02F_0|VDDR raven_padframe_0|FILLER02F_0|VDDO 0.06fF
C5763 BU_3VX2_8|A BU_3VX2_38|A 0.89fF
C5764 BU_3VX2_70|A BU_3VX2_64|A 1.94fF
C5765 BU_3VX2_17|A raven_soc_0|flash_clk 0.01fF
C5766 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_out<8> 0.43fF
C5767 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<9> 0.57fF
C5768 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<13> 0.18fF
C5769 raven_soc_0|gpio_in<0> BU_3VX2_29|Q 0.01fF
C5770 raven_soc_0|ram_wenb apllc03_1v8_0|CLK 0.47fF
C5771 raven_soc_0|gpio_out<13> BU_3VX2_27|Q 0.01fF
C5772 raven_soc_0|flash_csb BU_3VX2_29|Q 15.50fF
C5773 BU_3VX2_54|A BU_3VX2_55|Q 0.15fF
C5774 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<3> 1.02fF
C5775 BU_3VX2_9|A BU_3VX2_17|A 1.54fF
C5776 LS_3VX2_9|Q LS_3VX2_4|Q 6.72fF
C5777 raven_spi_0|SDI raven_soc_0|gpio_pullup<15> 1.48fF
C5778 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<15> 0.09fF
C5779 IN_3VX2_1|A raven_soc_0|gpio_pullup<7> 0.01fF
C5780 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<10> 0.01fF
C5781 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<5> 0.01fF
C5782 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<12> 10.93fF
C5783 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<10> 0.20fF
C5784 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_outenb<5> 0.03fF
C5785 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<15> 0.58fF
C5786 LS_3VX2_3|A raven_soc_0|gpio_out<11> 0.01fF
C5787 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<14> 0.02fF
C5788 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<9> 7.05fF
C5789 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<8> 0.56fF
C5790 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<18> 0.64fF
C5791 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<4> 0.17fF
C5792 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<7> 4.17fF
C5793 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<24> 0.21fF
C5794 AMUX4_3V_3|SEL[1] BU_3VX2_21|Q 1.55fF
C5795 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<22> 0.05fF
C5796 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<5> 2.98fF
C5797 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<25> 25.71fF
C5798 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<2> 0.17fF
C5799 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<12> 0.34fF
C5800 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<15> 13.74fF
C5801 AMUX4_3V_3|SEL[1] BU_3VX2_8|Q 0.01fF
C5802 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<8> 0.18fF
C5803 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<14> 0.02fF
C5804 raven_soc_0|ext_clk raven_soc_0|flash_io0_do 23.52fF
C5805 BU_3VX2_14|Q BU_3VX2_69|Q 4.09fF
C5806 BU_3VX2_70|Q BU_3VX2_68|Q 15.08fF
C5807 raven_soc_0|flash_io1_oeb VDD3V3 12.31fF
C5808 AMUX4_3V_4|AIN2 LS_3VX2_15|A 0.01fF
C5809 vdd BU_3VX2_24|Q 0.85fF
C5810 AMUX4_3V_0|SEL[0] BU_3VX2_72|Q 0.02fF
C5811 BU_3VX2_23|A BU_3VX2_35|A 0.01fF
C5812 raven_soc_0|gpio_pullup<2> BU_3VX2_63|Q 0.01fF
C5813 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<4> 10.54fF
C5814 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<6> 0.01fF
C5815 raven_padframe_0|aregc01_3v3_0|m4_92500_28769# raven_padframe_0|aregc01_3v3_0|GNDO 0.04fF
C5816 raven_padframe_0|aregc01_3v3_0|m4_0_22024# raven_padframe_0|aregc01_3v3_0|VDDO 1.17fF
C5817 AMUX4_3V_1|AIN1 BU_3VX2_59|A 0.02fF
C5818 BU_3VX2_68|A BU_3VX2_66|Q 0.03fF
C5819 BU_3VX2_12|A BU_3VX2_10|Q 0.03fF
C5820 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<31> 10.51fF
C5821 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<27> 0.11fF
C5822 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<25> 0.07fF
C5823 LS_3VX2_19|A BU_3VX2_60|Q 15.47fF
C5824 LS_3VX2_22|A BU_3VX2_58|Q 0.02fF
C5825 BU_3VX2_60|Q BU_3VX2_52|Q 16.84fF
C5826 BU_3VX2_24|A BU_3VX2_21|Q 0.02fF
C5827 BU_3VX2_2|A BU_3VX2_37|Q 0.16fF
C5828 AMUX4_3V_0|AIN1 LS_3VX2_27|Q 1.47fF
C5829 BU_3VX2_12|A raven_soc_0|flash_clk 0.01fF
C5830 BU_3VX2_13|A vdd 0.06fF
C5831 BU_3VX2_31|A apllc03_1v8_0|B_VCO 0.49fF
C5832 raven_soc_0|gpio_pulldown<14> raven_soc_0|ext_clk 0.01fF
C5833 BU_3VX2_0|Q LS_3VX2_18|A 10.23fF
C5834 raven_soc_0|gpio_pulldown<1> BU_3VX2_23|Q 0.01fF
C5835 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<5> 0.01fF
C5836 LS_3VX2_13|A VDD3V3 0.51fF
C5837 raven_soc_0|gpio_in<2> BU_3VX2_24|Q 0.48fF
C5838 raven_soc_0|gpio_outenb<13> BU_3VX2_71|Q 0.27fF
C5839 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<31> 0.01fF
C5840 BU_3VX2_11|Q BU_3VX2_36|Q 1.57fF
C5841 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<10> 0.02fF
C5842 raven_padframe_0|ICFC_1|GNDR raven_padframe_0|ICFC_1|VDDO 0.09fF
C5843 markings_0|manufacturer_0|_alphabet_F_0|m2_0_0# markings_0|manufacturer_0|_alphabet_E_1|m2_0_0# 0.38fF
C5844 markings_0|product_name_0|_alphabet_N_0|m2_0_0# markings_0|product_name_0|_alphabet_E_0|m2_0_0# 0.50fF
C5845 BU_3VX2_9|A BU_3VX2_12|A 4.56fF
C5846 BU_3VX2_66|A BU_3VX2_70|A 3.35fF
C5847 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_out<4> 0.51fF
C5848 raven_soc_0|gpio_pullup<0> BU_3VX2_0|Q 0.01fF
C5849 AMUX4_3V_4|AIN1 raven_soc_0|ser_rx 4.80fF
C5850 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<5> 0.01fF
C5851 raven_soc_0|gpio_in<0> raven_soc_0|flash_io2_do 0.13fF
C5852 raven_soc_0|gpio_in<3> raven_soc_0|flash_io1_di 2.33fF
C5853 BU_3VX2_36|A BU_3VX2_36|Q 0.08fF
C5854 raven_soc_0|gpio_in<4> apllc03_1v8_0|CLK 0.05fF
C5855 adc_low BU_3VX2_60|Q 0.05fF
C5856 raven_soc_0|flash_csb raven_soc_0|flash_io2_do 18.45fF
C5857 BU_3VX2_24|A BU_3VX2_19|A 4.39fF
C5858 raven_soc_0|gpio_in<9> raven_soc_0|irq_pin 0.01fF
C5859 BU_3VX2_73|Q BU_3VX2_49|Q 10.92fF
C5860 raven_soc_0|irq_pin BU_3VX2_42|Q 0.01fF
C5861 VDD raven_padframe_0|BBCUD4F_12|VDDR 0.71fF
C5862 LS_3VX2_12|Q LS_3VX2_11|Q 4.62fF
C5863 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<0> 138.34fF
C5864 BU_3VX2_17|A BU_3VX2_28|A 1.93fF
C5865 LS_3VX2_24|A LS_3VX2_24|Q 0.05fF
C5866 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_outenb<2> 32.70fF
C5867 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<10> 0.90fF
C5868 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<7> 9.38fF
C5869 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<6> 85.55fF
C5870 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<9> 0.01fF
C5871 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<8> 4.45fF
C5872 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<1> 10.93fF
C5873 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<17> 8.78fF
C5874 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<27> 3.16fF
C5875 BU_3VX2_1|Q BU_3VX2_7|Q 0.13fF
C5876 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<29> 0.01fF
C5877 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<19> 0.01fF
C5878 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<13> 0.01fF
C5879 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<26> 0.01fF
C5880 raven_soc_0|gpio_out<15> vdd 1.38fF
C5881 raven_soc_0|gpio_in<7> apllc03_1v8_0|CLK 0.02fF
C5882 AMUX4_3V_1|SEL[1] AMUX4_3V_4|AIN2 0.01fF
C5883 raven_soc_0|gpio_in<15> BU_3VX2_25|Q 0.01fF
C5884 raven_soc_0|gpio_in<11> BU_3VX2_24|Q 0.01fF
C5885 raven_soc_0|gpio_in<13> BU_3VX2_29|Q 0.01fF
C5886 raven_soc_0|gpio_in<14> BU_3VX2_27|Q 0.01fF
C5887 LS_3VX2_9|A LS_3VX2_12|A 14.68fF
C5888 raven_padframe_0|VDDPADFC_0|GNDR raven_padframe_0|VDDPADFC_0|GNDO 0.81fF
C5889 raven_padframe_0|BBCUD4F_12|VDDR LOGIC0_3V_4|Q 0.01fF
C5890 BU_3VX2_35|A IN_3VX2_1|A 0.01fF
C5891 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_out<2> 14.39fF
C5892 raven_padframe_0|aregc01_3v3_1|m4_92500_29333# raven_padframe_0|aregc01_3v3_1|m4_92500_28769# 0.03fF
C5893 IN_3VX2_1|A raven_soc_0|gpio_pulldown<15> 0.01fF
C5894 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<9> 0.01fF
C5895 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<12> 35.60fF
C5896 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<10> 0.01fF
C5897 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<11> 0.02fF
C5898 BU_3VX2_63|Q raven_soc_0|gpio_outenb<14> 0.01fF
C5899 LS_3VX2_14|A LS_3VX2_20|A 7.21fF
C5900 LS_3VX2_3|A raven_soc_0|gpio_in<12> 0.01fF
C5901 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<6> 0.01fF
C5902 raven_soc_0|gpio_pulldown<10> raven_soc_0|ext_clk 0.01fF
C5903 raven_soc_0|gpio_pulldown<13> VDD3V3 0.07fF
C5904 raven_soc_0|ser_rx VDD3V3 3.65fF
C5905 raven_soc_0|gpio_in<5> vdd 0.07fF
C5906 raven_soc_0|gpio_out<10> BU_3VX2_28|Q 0.01fF
C5907 raven_soc_0|gpio_pullup<14> BU_3VX2_26|Q 0.01fF
C5908 LS_3VX2_23|A vdd 1.53fF
C5909 BU_3VX2_14|Q BU_3VX2_29|Q 0.90fF
C5910 BU_3VX2_70|Q BU_3VX2_24|Q 1.75fF
C5911 BU_3VX2_37|Q apllc03_1v8_0|CLK 0.01fF
C5912 BU_3VX2_7|A raven_soc_0|flash_io0_di 0.01fF
C5913 BU_3VX2_20|A raven_soc_0|flash_io2_do 0.01fF
C5914 BU_3VX2_18|A raven_soc_0|flash_io2_oeb 0.01fF
C5915 raven_padframe_0|BT4F_2|VDDR raven_padframe_0|BT4F_2|GNDO 0.13fF
C5916 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<15> 3.82fF
C5917 BU_3VX2_31|A raven_soc_0|flash_io3_do 4.68fF
C5918 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<10> 5.31fF
C5919 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<3> 3.74fF
C5920 BU_3VX2_0|Q raven_soc_0|ram_wdata<31> 0.02fF
C5921 raven_soc_0|gpio_pullup<1> VDD3V3 1.97fF
C5922 VDD raven_padframe_0|axtoc02_3v3_0|m4_55000_31172# 0.25fF
C5923 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<0> 1.04fF
C5924 BU_3VX2_48|A BU_3VX2_47|A 10.09fF
C5925 BU_3VX2_51|A BU_3VX2_45|A 0.50fF
C5926 BU_3VX2_60|Q BU_3VX2_58|Q 81.21fF
C5927 BU_3VX2_41|A adc0_data<5> 0.10fF
C5928 raven_padframe_0|BBCUD4F_11|GNDR raven_padframe_0|BBCUD4F_11|GNDO 0.81fF
C5929 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<0> 30.66fF
C5930 BU_3VX2_6|A BU_3VX2_18|A 0.91fF
C5931 BU_3VX2_68|A BU_3VX2_0|Q 1.11fF
C5932 BU_3VX2_12|A BU_3VX2_28|A 0.01fF
C5933 BU_3VX2_23|A raven_soc_0|flash_io3_di 0.01fF
C5934 raven_soc_0|gpio_out<0> BU_3VX2_23|Q 0.01fF
C5935 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<13> 0.12fF
C5936 BU_3VX2_31|A raven_soc_0|gpio_out<14> 0.01fF
C5937 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<5> 0.49fF
C5938 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<6> 0.01fF
C5939 raven_soc_0|gpio_out<13> BU_3VX2_25|Q 0.01fF
C5940 raven_soc_0|gpio_out<7> apllc03_1v8_0|CLK 0.01fF
C5941 raven_soc_0|gpio_out<12> BU_3VX2_23|Q 0.01fF
C5942 raven_soc_0|gpio_outenb<15> BU_3VX2_27|Q 0.01fF
C5943 raven_soc_0|gpio_out<9> BU_3VX2_28|Q 0.01fF
C5944 BU_3VX2_54|A BU_3VX2_57|Q 0.02fF
C5945 BU_3VX2_56|Q LS_3VX2_20|A 0.10fF
C5946 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<5> 0.01fF
C5947 BU_3VX2_19|A BU_3VX2_16|A 7.19fF
C5948 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<4> 0.31fF
C5949 BU_3VX2_19|A BU_3VX2_29|A 2.09fF
C5950 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<6> 0.01fF
C5951 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<12> 0.01fF
C5952 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<15> 0.02fF
C5953 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<10> 0.27fF
C5954 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<7> 2.70fF
C5955 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<5> 2.43fF
C5956 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<9> 0.01fF
C5957 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<10> 45.08fF
C5958 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<8> 0.01fF
C5959 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<9> 0.01fF
C5960 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<7> 4.73fF
C5961 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<20> 0.01fF
C5962 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<10> 79.44fF
C5963 AMUX4_3V_3|SEL[1] BU_3VX2_19|Q 0.01fF
C5964 raven_spi_0|CSB raven_spi_0|SDI 70.88fF
C5965 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<12> 6.93fF
C5966 AMUX4_3V_3|SEL[1] BU_3VX2_18|Q 0.71fF
C5967 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<0> 1.40fF
C5968 raven_soc_0|gpio_in<11> raven_soc_0|gpio_out<15> 1.85fF
C5969 BU_3VX2_40|Q raven_soc_0|flash_io3_oeb 0.01fF
C5970 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<1> 2.29fF
C5971 raven_soc_0|ext_clk raven_soc_0|flash_io1_di 85.38fF
C5972 raven_padframe_0|FILLER20F_8|GNDR raven_padframe_0|FILLER20F_8|GNDO 0.81fF
C5973 BU_3VX2_17|A BU_3VX2_14|A 8.06fF
C5974 IN_3VX2_1|A raven_soc_0|gpio_pulldown<0> 0.01fF
C5975 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<8> 0.01fF
C5976 raven_padframe_0|aregc01_3v3_0|m4_92500_29057# raven_padframe_0|aregc01_3v3_0|m4_92500_28769# 0.11fF
C5977 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<14> 0.48fF
C5978 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_outenb<6> 0.30fF
C5979 AMUX4_3V_1|AIN1 AMUX4_3V_1|AOUT 0.80fF
C5980 adc_high raven_soc_0|irq_pin 0.25fF
C5981 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<28> 5.52fF
C5982 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<11> 1.20fF
C5983 BU_3VX2_71|Q raven_soc_0|gpio_in<8> 0.10fF
C5984 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<11> 0.32fF
C5985 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<19> 12.26fF
C5986 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<23> 0.04fF
C5987 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_out<15> 0.02fF
C5988 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<7> 7.80fF
C5989 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<17> 0.02fF
C5990 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<19> 0.01fF
C5991 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<14> 0.03fF
C5992 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<2> 11.27fF
C5993 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<26> 0.02fF
C5994 LS_3VX2_19|A BU_3VX2_62|Q 33.87fF
C5995 raven_soc_0|ram_wdata<20> vdd 0.86fF
C5996 LS_3VX2_22|A BU_3VX2_60|Q 0.02fF
C5997 BU_3VX2_62|Q BU_3VX2_52|Q 13.37fF
C5998 BU_3VX2_35|A BU_3VX2_25|A 0.01fF
C5999 raven_padframe_0|POWERCUTVDD3FC_1|VDDR LOGIC0_3V_4|Q 0.01fF
C6000 acsoc02_3v3_0|CS_8U VDD3V3 0.02fF
C6001 IN_3VX2_1|A BU_3VX2_30|Q 0.08fF
C6002 raven_soc_0|gpio_outenb<4> BU_3VX2_40|Q 0.17fF
C6003 LS_3VX2_5|A LS_3VX2_19|A 0.01fF
C6004 LS_3VX2_5|A BU_3VX2_52|Q 18.50fF
C6005 BU_3VX2_69|A BU_3VX2_68|Q 0.16fF
C6006 raven_soc_0|gpio_outenb<1> BU_3VX2_29|Q 0.01fF
C6007 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_outenb<13> 14.74fF
C6008 raven_soc_0|gpio_out<8> raven_soc_0|gpio_out<14> 1.22fF
C6009 raven_soc_0|gpio_pullup<13> BU_3VX2_71|Q 0.13fF
C6010 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<5> 0.01fF
C6011 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<31> 2.57fF
C6012 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<10> 4.19fF
C6013 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<9> 0.10fF
C6014 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<6> 0.74fF
C6015 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<24> 0.01fF
C6016 raven_padframe_0|ICF_2|GNDR raven_padframe_0|ICF_2|VDDO 0.09fF
C6017 markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# markings_0|manufacturer_0|_alphabet_F_0|m2_0_0# 0.02fF
C6018 BU_3VX2_3|A raven_soc_0|flash_io3_oeb 0.01fF
C6019 BU_3VX2_22|A raven_soc_0|flash_io3_do 0.01fF
C6020 AMUX4_3V_3|AOUT raven_soc_0|flash_io1_do 1.66fF
C6021 BU_3VX2_15|A raven_soc_0|flash_io3_oeb 0.01fF
C6022 raven_soc_0|gpio_pullup<2> BU_3VX2_24|Q 0.01fF
C6023 BU_3VX2_71|A raven_soc_0|flash_io2_oeb 0.01fF
C6024 VDD raven_padframe_0|FILLER20F_0|GNDO 0.07fF
C6025 IN_3VX2_1|A raven_soc_0|flash_io3_di 3.80fF
C6026 VDD raven_padframe_0|VDDORPADF_0|GNDR 0.16fF
C6027 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<10> 27.10fF
C6028 adc_low BU_3VX2_62|Q 0.05fF
C6029 BU_3VX2_3|A BU_3VX2_2|A 16.39fF
C6030 BU_3VX2_7|A BU_3VX2_5|A 8.95fF
C6031 BU_3VX2_23|A BU_3VX2_63|A 0.01fF
C6032 BU_3VX2_6|A BU_3VX2_71|A 0.02fF
C6033 BU_3VX2_19|A LS_3VX2_3|Q 0.01fF
C6034 BU_3VX2_2|A BU_3VX2_15|A 0.97fF
C6035 BU_3VX2_8|A BU_3VX2_31|A 0.01fF
C6036 BU_3VX2_31|A raven_soc_0|gpio_pulldown<1> 0.01fF
C6037 BU_3VX2_18|A BU_3VX2_27|A 2.39fF
C6038 BU_3VX2_12|A BU_3VX2_14|A 11.89fF
C6039 AMUX4_3V_0|AIN1 BU_3VX2_41|A 0.02fF
C6040 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<14> 0.16fF
C6041 raven_soc_0|gpio_out<5> BU_3VX2_71|Q 0.01fF
C6042 raven_soc_0|gpio_out<7> raven_soc_0|gpio_outenb<8> 4.81fF
C6043 AMUX2_3V_0|SEL BU_3VX2_59|Q 0.13fF
C6044 BU_3VX2_13|Q BU_3VX2_66|Q 1.02fF
C6045 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<29> 63.11fF
C6046 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<2> 0.17fF
C6047 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<21> 0.01fF
C6048 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<7> 0.01fF
C6049 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<27> 6.61fF
C6050 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<6> 0.01fF
C6051 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<25> 0.01fF
C6052 BU_3VX2_2|Q BU_3VX2_10|Q 26.00fF
C6053 BU_3VX2_21|Q BU_3VX2_67|Q 6.43fF
C6054 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<1> 1.32fF
C6055 BU_3VX2_13|Q BU_3VX2_20|Q 4.73fF
C6056 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<26> 2.98fF
C6057 BU_3VX2_38|Q BU_3VX2_8|Q 4.92fF
C6058 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<21> 7.98fF
C6059 LS_3VX2_18|A AMUX4_3V_3|SEL[0] 1.01fF
C6060 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<25> 5.54fF
C6061 BU_3VX2_67|Q BU_3VX2_8|Q 8.09fF
C6062 BU_3VX2_40|Q apllc03_1v8_0|CLK 89.65fF
C6063 raven_soc_0|gpio_in<6> vdd 1.57fF
C6064 BU_3VX2_22|Q BU_3VX2_17|Q 6.93fF
C6065 raven_soc_0|ext_clk BU_3VX2_28|Q 0.01fF
C6066 raven_soc_0|gpio_in<9> BU_3VX2_26|Q 0.01fF
C6067 raven_soc_0|gpio_in<14> BU_3VX2_25|Q 0.01fF
C6068 AMUX4_3V_0|SEL[1] BU_3VX2_43|Q 163.64fF
C6069 BU_3VX2_43|Q BU_3VX2_51|Q 12.91fF
C6070 BU_3VX2_55|Q BU_3VX2_53|Q 80.18fF
C6071 LS_3VX2_15|Q vdd 0.48fF
C6072 raven_padframe_0|APR00DF_2|GNDR raven_padframe_0|APR00DF_2|VDDO 0.09fF
C6073 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<7> 0.64fF
C6074 raven_padframe_0|axtoc02_3v3_0|m4_0_30133# raven_padframe_0|axtoc02_3v3_0|m4_0_29057# 0.02fF
C6075 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<9> 0.01fF
C6076 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<3> 0.01fF
C6077 BU_3VX2_63|Q raven_soc_0|gpio_pullup<15> 0.01fF
C6078 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<10> 0.01fF
C6079 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<12> 16.93fF
C6080 BU_3VX2_10|A raven_soc_0|ext_clk 0.08fF
C6081 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<5> 0.73fF
C6082 raven_soc_0|gpio_pulldown<12> raven_soc_0|ext_clk 0.01fF
C6083 raven_soc_0|gpio_out<10> vdd 0.21fF
C6084 AMUX4_3V_3|SEL[1] BU_3VX2_27|Q 0.07fF
C6085 BU_3VX2_56|Q BU_3VX2_47|Q 1.32fF
C6086 raven_soc_0|gpio_in<6> raven_padframe_0|BBCUD4F_6|PO 0.04fF
C6087 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<11> 1.81fF
C6088 BU_3VX2_9|A BU_3VX2_10|Q 0.03fF
C6089 VDD raven_padframe_0|FILLER50F_2|GNDR 0.16fF
C6090 BU_3VX2_0|A raven_soc_0|ext_clk 79.94fF
C6091 IN_3VX2_1|Q AMUX4_3V_4|AIN2 4.09fF
C6092 VDD raven_padframe_0|FILLER20F_7|GNDR 0.16fF
C6093 IN_3VX2_1|A raven_soc_0|irq_pin 95.89fF
C6094 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<6> 0.47fF
C6095 LS_3VX2_5|Q vdd 0.09fF
C6096 VDD raven_padframe_0|BBCUD4F_10|GNDO 0.07fF
C6097 LS_3VX2_3|A raven_soc_0|gpio_pulldown<7> 0.72fF
C6098 BU_3VX2_0|Q raven_soc_0|ram_wdata<19> 0.02fF
C6099 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<16> 0.31fF
C6100 BU_3VX2_51|A BU_3VX2_50|A 13.29fF
C6101 BU_3VX2_62|Q BU_3VX2_58|Q 29.26fF
C6102 BU_3VX2_61|Q BU_3VX2_59|Q 81.44fF
C6103 raven_padframe_0|BBCUD4F_4|VDDO raven_padframe_0|BBCUD4F_4|GNDO 2.28fF
C6104 raven_soc_0|gpio_in<1> BU_3VX2_29|Q 0.01fF
C6105 BU_3VX2_21|A raven_soc_0|flash_io3_do 0.10fF
C6106 BU_3VX2_9|A raven_soc_0|flash_clk 0.01fF
C6107 BU_3VX2_19|A raven_soc_0|flash_io1_oeb 0.01fF
C6108 BU_3VX2_17|A raven_soc_0|flash_io1_do 0.01fF
C6109 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<13> 0.29fF
C6110 raven_padframe_0|ICFC_2|VDDR raven_padframe_0|ICFC_2|GNDR 0.68fF
C6111 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<15> 3.07fF
C6112 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<10> 0.01fF
C6113 LS_3VX2_5|A BU_3VX2_58|Q 8.46fF
C6114 raven_soc_0|gpio_in<3> vdd 2.32fF
C6115 VDD raven_padframe_0|FILLER10F_0|GNDR 0.16fF
C6116 raven_soc_0|gpio_out<9> vdd 0.23fF
C6117 raven_soc_0|gpio_outenb<7> apllc03_1v8_0|CLK 0.01fF
C6118 raven_soc_0|gpio_outenb<12> BU_3VX2_23|Q 0.01fF
C6119 raven_soc_0|gpio_outenb<15> BU_3VX2_25|Q 0.01fF
C6120 raven_soc_0|gpio_outenb<10> BU_3VX2_28|Q 0.01fF
C6121 raven_soc_0|gpio_outenb<14> BU_3VX2_24|Q 0.01fF
C6122 LS_3VX2_12|Q LS_3VX2_8|A 0.54fF
C6123 BU_3VX2_63|A IN_3VX2_1|A 0.01fF
C6124 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<12> 0.17fF
C6125 BU_3VX2_0|Q raven_soc_0|gpio_pullup<3> 0.01fF
C6126 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<10> 6.08fF
C6127 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<10> 146.45fF
C6128 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<7> 1.37fF
C6129 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_outenb<0> 0.01fF
C6130 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<8> 0.01fF
C6131 BU_3VX2_25|A raven_soc_0|flash_io3_di 0.01fF
C6132 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<14> 0.10fF
C6133 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<4> 0.02fF
C6134 raven_soc_0|gpio_in<6> raven_soc_0|gpio_in<11> 24.96fF
C6135 raven_soc_0|gpio_in<7> raven_soc_0|gpio_in<15> 16.91fF
C6136 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<10> 12.52fF
C6137 AMUX4_3V_3|SEL[1] AMUX4_3V_4|SEL[1] 34.14fF
C6138 LS_3VX2_16|Q LS_3VX2_17|Q 13.70fF
C6139 LS_3VX2_15|Q BU_3VX2_62|A 2.05fF
C6140 VDD3V3 AMUX4_3V_1|SEL[0] 0.71fF
C6141 AMUX4_3V_0|SEL[1] BU_3VX2_50|Q 10.29fF
C6142 BU_3VX2_22|A BU_3VX2_8|A 0.68fF
C6143 VDD raven_padframe_0|ICF_0|VDDR 0.71fF
C6144 BU_3VX2_50|Q BU_3VX2_51|Q 211.84fF
C6145 raven_padframe_0|BT4F_2|GNDR raven_padframe_0|BT4F_2|VDDO 0.09fF
C6146 BU_3VX2_35|A BU_3VX2_4|A 1.51fF
C6147 raven_soc_0|gpio_out<0> BU_3VX2_31|A 0.01fF
C6148 BU_3VX2_0|A BU_3VX2_65|A 1.51fF
C6149 BU_3VX2_71|A BU_3VX2_27|A 0.01fF
C6150 raven_padframe_0|APR00DF_0|GNDR raven_padframe_0|APR00DF_0|GNDO 0.81fF
C6151 raven_padframe_0|FILLER20F_4|VDDO raven_padframe_0|FILLER20F_4|GNDO 2.28fF
C6152 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<3> 7.81fF
C6153 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<3> 0.55fF
C6154 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<9> 0.01fF
C6155 BU_3VX2_31|A raven_soc_0|gpio_out<12> 0.01fF
C6156 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<8> 0.10fF
C6157 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<15> 0.21fF
C6158 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<11> 0.02fF
C6159 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<8> 0.01fF
C6160 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<28> 2.19fF
C6161 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<11> 10.31fF
C6162 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<20> 0.01fF
C6163 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<0> 0.31fF
C6164 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<19> 0.21fF
C6165 raven_soc_0|gpio_outenb<8> BU_3VX2_40|Q 0.01fF
C6166 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<11> 0.01fF
C6167 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<6> 0.01fF
C6168 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<9> 0.01fF
C6169 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<2> 0.02fF
C6170 LS_3VX2_22|A BU_3VX2_62|Q 0.02fF
C6171 BU_3VX2_71|Q VDD3V3 0.67fF
C6172 raven_soc_0|ram_rdata<21> vdd 0.36fF
C6173 raven_padframe_0|ICF_0|VDDR LOGIC0_3V_4|Q 0.01fF
C6174 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<1> 135.13fF
C6175 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<13> 0.67fF
C6176 raven_soc_0|gpio_out<3> BU_3VX2_63|Q 0.01fF
C6177 LS_3VX2_2|Q VDD3V3 0.26fF
C6178 LS_3VX2_5|A LS_3VX2_22|A 8.80fF
C6179 BU_3VX2_12|A raven_soc_0|flash_io1_do 0.01fF
C6180 BU_3VX2_0|Q BU_3VX2_13|Q 0.01fF
C6181 raven_soc_0|gpio_pullup<0> BU_3VX2_26|Q 0.01fF
C6182 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<30> 9.17fF
C6183 raven_soc_0|ram_rdata<14> raven_soc_0|ram_addr<2> 0.01fF
C6184 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<6> 10.51fF
C6185 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_pullup<14> 32.69fF
C6186 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<9> 4.51fF
C6187 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<24> 0.02fF
C6188 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<31> 9.06fF
C6189 raven_soc_0|gpio_out<10> raven_soc_0|gpio_outenb<9> 15.80fF
C6190 raven_soc_0|ram_rdata<4> raven_soc_0|ram_addr<4> 0.13fF
C6191 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<7> 0.01fF
C6192 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_out<14> 0.02fF
C6193 raven_soc_0|ram_wdata<23> raven_soc_0|ram_addr<3> 0.01fF
C6194 BU_3VX2_14|Q BU_3VX2_32|Q 2.93fF
C6195 raven_padframe_0|APR00DF_1|GNDR raven_padframe_0|APR00DF_1|GNDO 0.81fF
C6196 raven_padframe_0|axtoc02_3v3_0|VDDR raven_padframe_0|axtoc02_3v3_0|GNDO 0.19fF
C6197 BU_3VX2_24|A raven_soc_0|flash_io2_oeb 2.98fF
C6198 raven_padframe_0|GNDORPADF_5|VDDR raven_padframe_0|GNDORPADF_5|VDDO 0.06fF
C6199 VDD raven_padframe_0|GNDORPADF_5|GNDOR 0.24fF
C6200 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<12> 0.03fF
C6201 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<11> 0.06fF
C6202 VDD raven_padframe_0|GNDORPADF_0|VDDR 0.71fF
C6203 BU_3VX2_28|A raven_soc_0|flash_clk 9.90fF
C6204 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<13> 6.86fF
C6205 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<15> 0.16fF
C6206 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<7> 0.22fF
C6207 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<11> 4.78fF
C6208 BU_3VX2_29|A BU_3VX2_27|Q 0.03fF
C6209 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<15> 33.73fF
C6210 VDD raven_padframe_0|VDDORPADF_1|GNDR 0.16fF
C6211 raven_padframe_0|APR00DF_1|VDDR raven_padframe_0|APR00DF_1|GNDO 0.13fF
C6212 BU_3VX2_24|A BU_3VX2_6|A 0.01fF
C6213 raven_spi_0|SDI BU_3VX2_2|A 0.01fF
C6214 BU_3VX2_9|A BU_3VX2_28|A 0.01fF
C6215 BU_3VX2_7|A BU_3VX2_13|A 1.96fF
C6216 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<2> 13.05fF
C6217 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<8> 0.28fF
C6218 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<9> 0.01fF
C6219 raven_soc_0|gpio_outenb<6> BU_3VX2_71|Q 0.01fF
C6220 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<14> 0.50fF
C6221 raven_soc_0|gpio_out<9> raven_soc_0|gpio_outenb<9> 96.96fF
C6222 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<8> 0.69fF
C6223 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<8> 10.23fF
C6224 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<5> 0.01fF
C6225 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pullup<14> 0.01fF
C6226 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<15> 0.01fF
C6227 AMUX2_3V_0|SEL BU_3VX2_61|Q 0.01fF
C6228 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_4|PO 0.04fF
C6229 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<2> 4.17fF
C6230 BU_3VX2_6|Q BU_3VX2_12|Q 6.26fF
C6231 BU_3VX2_19|Q BU_3VX2_38|Q 0.39fF
C6232 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<15> 0.48fF
C6233 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<17> 136.25fF
C6234 BU_3VX2_16|Q BU_3VX2_13|Q 13.52fF
C6235 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<14> 0.02fF
C6236 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<25> 58.76fF
C6237 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<21> 4.53fF
C6238 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<26> 7.33fF
C6239 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<1> 0.01fF
C6240 BU_3VX2_21|Q BU_3VX2_65|Q 22.62fF
C6241 BU_3VX2_13|Q BU_3VX2_30|Q 0.18fF
C6242 BU_3VX2_12|Q BU_3VX2_7|Q 10.84fF
C6243 BU_3VX2_18|Q BU_3VX2_67|Q 7.94fF
C6244 BU_3VX2_66|Q BU_3VX2_69|Q 9.67fF
C6245 BU_3VX2_19|Q BU_3VX2_67|Q 5.04fF
C6246 BU_3VX2_69|Q BU_3VX2_20|Q 0.01fF
C6247 BU_3VX2_38|Q BU_3VX2_18|Q 0.17fF
C6248 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<13> 35.76fF
C6249 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<17> 4.48fF
C6250 BU_3VX2_15|Q BU_3VX2_9|Q 6.04fF
C6251 raven_soc_0|ext_clk vdd 1.88fF
C6252 VDD3V3 LS_3VX2_17|A 0.92fF
C6253 BU_3VX2_43|Q BU_3VX2_49|Q 17.29fF
C6254 BU_3VX2_57|Q BU_3VX2_53|Q 34.66fF
C6255 BU_3VX2_52|A vdd 0.07fF
C6256 BU_3VX2_44|A BU_3VX2_44|Q 0.10fF
C6257 AMUX4_3V_0|SEL[0] BU_3VX2_42|Q 6.74fF
C6258 BU_3VX2_8|A BU_3VX2_21|A 1.17fF
C6259 raven_padframe_0|POWERCUTVDD3FC_1|GNDR raven_padframe_0|POWERCUTVDD3FC_1|GNDO 0.77fF
C6260 LOGIC1_3V_3|Q LOGIC0_3V_4|Q 2.90fF
C6261 BU_3VX2_25|A BU_3VX2_63|A 0.01fF
C6262 raven_padframe_0|BBCUD4F_10|GNDR raven_padframe_0|BBCUD4F_10|GNDO 0.81fF
C6263 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<9> 0.01fF
C6264 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<5> 0.19fF
C6265 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<4> 0.01fF
C6266 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<0> 0.01fF
C6267 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<3> 0.87fF
C6268 raven_soc_0|flash_clk BU_3VX2_33|Q 0.01fF
C6269 raven_soc_0|ram_rdata<17> vdd 0.38fF
C6270 AMUX4_3V_3|SEL[1] BU_3VX2_25|Q 0.88fF
C6271 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<6> 0.27fF
C6272 AMUX4_3V_3|AOUT raven_soc_0|flash_csb 9.16fF
C6273 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<2> 6.97fF
C6274 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<13> 0.47fF
C6275 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<12> 1.14fF
C6276 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<8> 0.03fF
C6277 VDD raven_padframe_0|FILLER40F_0|GNDO 0.07fF
C6278 VDD raven_padframe_0|FILLER20F_1|GNDR 0.16fF
C6279 BU_3VX2_40|A raven_soc_0|ext_clk 3.12fF
C6280 VDD raven_padframe_0|CORNERESDF_2|GNDO 0.07fF
C6281 raven_soc_0|gpio_in<2> raven_soc_0|ext_clk 0.01fF
C6282 BU_3VX2_0|Q raven_soc_0|ram_wdata<30> 0.02fF
C6283 raven_soc_0|gpio_outenb<3> VDD3V3 0.40fF
C6284 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<13> 0.08fF
C6285 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<15> 0.02fF
C6286 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<17> 3.13fF
C6287 raven_soc_0|flash_io2_di raven_soc_0|flash_io0_do 53.85fF
C6288 raven_soc_0|ram_addr<2> raven_soc_0|ram_addr<0> 33.05fF
C6289 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<1> 2.23fF
C6290 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<31> 3.59fF
C6291 LS_3VX2_2|A LS_3VX2_23|A 0.48fF
C6292 BU_3VX2_62|Q BU_3VX2_60|Q 58.54fF
C6293 LS_3VX2_15|A BU_3VX2_59|Q 36.14fF
C6294 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<1> 47.54fF
C6295 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<5> 0.96fF
C6296 raven_padframe_0|FILLER20F_3|VDDO raven_padframe_0|FILLER20F_3|GNDO 2.28fF
C6297 BU_3VX2_24|A BU_3VX2_25|Q 0.03fF
C6298 LS_3VX2_12|A BU_3VX2_73|Q 12.39fF
C6299 LS_3VX2_23|Q VDD3V3 0.46fF
C6300 BU_3VX2_16|A raven_soc_0|flash_io2_oeb 0.01fF
C6301 VDD BU_3VX2_27|Q 0.02fF
C6302 BU_3VX2_4|A raven_soc_0|flash_io3_di 0.06fF
C6303 LS_3VX2_11|A LS_3VX2_19|A 0.01fF
C6304 LS_3VX2_11|A BU_3VX2_52|Q 10.68fF
C6305 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<6> 0.93fF
C6306 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<14> 2.63fF
C6307 raven_padframe_0|ICF_2|VDDR raven_padframe_0|ICF_2|GNDO 0.13fF
C6308 BU_3VX2_29|A raven_soc_0|flash_io2_oeb 6.81fF
C6309 BU_3VX2_65|A vdd 0.22fF
C6310 IN_3VX2_1|A BU_3VX2_26|Q 34.55fF
C6311 LS_3VX2_5|A BU_3VX2_60|Q 6.47fF
C6312 raven_soc_0|gpio_outenb<10> vdd 0.26fF
C6313 VDD raven_padframe_0|FILLER20F_5|GNDR 0.16fF
C6314 raven_soc_0|gpio_pullup<12> BU_3VX2_23|Q 0.01fF
C6315 raven_soc_0|gpio_pullup<9> apllc03_1v8_0|CLK 0.01fF
C6316 raven_soc_0|gpio_pullup<15> BU_3VX2_24|Q 0.01fF
C6317 raven_soc_0|gpio_pullup<7> BU_3VX2_29|Q 0.01fF
C6318 raven_soc_0|gpio_pullup<10> BU_3VX2_28|Q 0.01fF
C6319 BU_3VX2_6|A BU_3VX2_16|A 1.10fF
C6320 BU_3VX2_6|A BU_3VX2_29|A 0.01fF
C6321 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<12> 0.01fF
C6322 BU_3VX2_37|A raven_soc_0|flash_io2_oeb 0.01fF
C6323 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<4> 0.36fF
C6324 LS_3VX2_3|A raven_soc_0|gpio_pullup<4> 0.01fF
C6325 BU_3VX2_35|A raven_soc_0|flash_io0_oeb 0.01fF
C6326 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<10> 9.52fF
C6327 raven_soc_0|gpio_pulldown<5> BU_3VX2_0|Q 0.01fF
C6328 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<6> 0.91fF
C6329 BU_3VX2_14|A raven_soc_0|flash_clk 0.01fF
C6330 LOGIC0_3V_4|Q BU_3VX2_27|Q 0.01fF
C6331 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<8> 25.02fF
C6332 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<13> 35.49fF
C6333 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<7> 0.43fF
C6334 raven_soc_0|ext_clk raven_soc_0|gpio_in<11> 0.01fF
C6335 BU_3VX2_40|Q raven_soc_0|gpio_in<15> 0.01fF
C6336 BU_3VX2_52|A BU_3VX2_62|A 0.12fF
C6337 BU_3VX2_56|A BU_3VX2_61|A 0.47fF
C6338 BU_3VX2_57|A BU_3VX2_60|A 1.06fF
C6339 BU_3VX2_58|A BU_3VX2_59|A 6.93fF
C6340 BU_3VX2_54|A LS_3VX2_16|Q 0.13fF
C6341 BU_3VX2_55|A LS_3VX2_15|Q 0.19fF
C6342 BU_3VX2_53|A LS_3VX2_17|Q 0.10fF
C6343 raven_soc_0|irq_pin BU_3VX2_54|Q 0.01fF
C6344 AMUX4_3V_0|SEL[1] BU_3VX2_48|Q 13.35fF
C6345 BU_3VX2_48|Q BU_3VX2_51|Q 50.65fF
C6346 BU_3VX2_49|Q BU_3VX2_50|Q 216.39fF
C6347 BU_3VX2_44|A vdd 0.06fF
C6348 BU_3VX2_24|A BU_3VX2_27|A 13.52fF
C6349 BU_3VX2_6|A BU_3VX2_37|A 1.68fF
C6350 LS_3VX2_13|Q LS_3VX2_10|Q 1.02fF
C6351 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<2> 3.92fF
C6352 BU_3VX2_9|A BU_3VX2_14|A 2.56fF
C6353 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<5> 3.17fF
C6354 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<6> 1.44fF
C6355 BU_3VX2_31|A raven_soc_0|gpio_outenb<12> 0.01fF
C6356 raven_padframe_0|aregc01_3v3_0|m4_0_31172# raven_padframe_0|aregc01_3v3_0|m4_0_30653# 0.09fF
C6357 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<10> 0.01fF
C6358 markings_0|efabless_logo_0|m1_0_n4950# markings_0|efabless_logo_0|m1_1500_n9450# 0.36fF
C6359 markings_0|efabless_logo_0|m1_8700_n6150# markings_0|efabless_logo_0|m1_8400_n7350# 0.28fF
C6360 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<10> 0.02fF
C6361 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<7> 7.28fF
C6362 raven_soc_0|gpio_outenb<9> raven_soc_0|ext_clk 0.01fF
C6363 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<9> 0.01fF
C6364 raven_soc_0|gpio_out<8> raven_soc_0|gpio_pullup<5> 0.80fF
C6365 raven_soc_0|gpio_pullup<14> VDD3V3 0.07fF
C6366 LS_3VX2_16|A BU_3VX2_53|Q 8.56fF
C6367 BU_3VX2_66|Q BU_3VX2_29|Q 0.01fF
C6368 BU_3VX2_20|Q BU_3VX2_29|Q 13.48fF
C6369 BU_3VX2_67|Q BU_3VX2_27|Q 3.62fF
C6370 BU_3VX2_38|Q BU_3VX2_27|Q 1.71fF
C6371 BU_3VX2_17|Q apllc03_1v8_0|CLK 0.01fF
C6372 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_in<3> 6.19fF
C6373 BU_3VX2_17|A raven_soc_0|flash_csb 0.01fF
C6374 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<15> 0.01fF
C6375 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<14> 1.56fF
C6376 LS_3VX2_12|Q vdd 0.97fF
C6377 LS_3VX2_24|A BU_3VX2_51|Q 9.07fF
C6378 VDD raven_padframe_0|APR00DF_3|VDDR 0.71fF
C6379 BU_3VX2_0|Q BU_3VX2_69|Q 0.01fF
C6380 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<24> 37.14fF
C6381 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<23> 3.30fF
C6382 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<14> 15.50fF
C6383 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<8> 57.40fF
C6384 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<30> 10.38fF
C6385 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<4> 45.57fF
C6386 AMUX4_3V_1|SEL[1] BU_3VX2_59|Q 11.06fF
C6387 raven_soc_0|flash_io1_oeb BU_3VX2_27|Q 0.01fF
C6388 adc0_data<5> BU_3VX2_72|Q 1.45fF
C6389 raven_padframe_0|axtoc02_3v3_0|m4_55000_22024# raven_padframe_0|axtoc02_3v3_0|VDDO 2.34fF
C6390 markings_0|mask_copyright_0|m2_n208_960# markings_0|manufacturer_0|_alphabet_E_1|m2_0_0# 0.03fF
C6391 markings_0|manufacturer_0|_alphabet_S_0|m2_32_224# markings_0|product_name_0|_alphabet_V_1|m2_0_560# 0.16fF
C6392 LS_3VX2_3|Q raven_soc_0|flash_io2_oeb 0.01fF
C6393 LS_3VX2_7|A BU_3VX2_59|Q 0.01fF
C6394 VDD raven_padframe_0|BBCUD4F_12|GNDR 0.16fF
C6395 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<7> 0.70fF
C6396 AMUX2_3V_0|AOUT AMUX4_3V_4|AIN3 0.68fF
C6397 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<14> 0.03fF
C6398 LS_3VX2_6|A BU_3VX2_54|Q 10.07fF
C6399 raven_soc_0|gpio_out<13> BU_3VX2_40|Q 0.05fF
C6400 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<9> 0.62fF
C6401 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<6> 0.12fF
C6402 LS_3VX2_3|A raven_soc_0|flash_clk 0.58fF
C6403 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<15> 0.02fF
C6404 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<11> 11.72fF
C6405 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pullup<5> 15.50fF
C6406 BU_3VX2_0|Q raven_soc_0|flash_io0_oeb 0.01fF
C6407 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<15> 48.78fF
C6408 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<23> 10.68fF
C6409 BU_3VX2_6|A LS_3VX2_3|Q 0.53fF
C6410 VDD raven_padframe_0|BBCUD4F_7|VDDR 0.71fF
C6411 BU_3VX2_63|A BU_3VX2_4|A 0.01fF
C6412 BU_3VX2_68|A BU_3VX2_36|A 2.45fF
C6413 analog_out adc_high 5.38fF
C6414 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<6> 0.01fF
C6415 LOGIC0_3V_4|Q raven_soc_0|flash_io2_oeb 0.01fF
C6416 BU_3VX2_25|A BU_3VX2_26|Q 0.03fF
C6417 IN_3VX2_1|A raven_soc_0|gpio_outenb<13> 0.01fF
C6418 LS_3VX2_11|A BU_3VX2_58|Q 0.01fF
C6419 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<7> 0.01fF
C6420 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<8> 0.02fF
C6421 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pullup<14> 1.36fF
C6422 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<10> 0.30fF
C6423 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<9> 15.03fF
C6424 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<5> 0.01fF
C6425 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<14> 8.34fF
C6426 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pullup<6> 39.39fF
C6427 raven_soc_0|gpio_pullup<8> BU_3VX2_71|Q 0.01fF
C6428 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<8> 5.77fF
C6429 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pulldown<6> 0.02fF
C6430 raven_padframe_0|BBCUD4F_9|VDDR raven_padframe_0|BBCUD4F_9|GNDR 0.68fF
C6431 AMUX2_3V_0|SEL LS_3VX2_15|A 0.02fF
C6432 raven_soc_0|gpio_pulldown<15> BU_3VX2_29|Q 0.01fF
C6433 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<3> 0.20fF
C6434 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<28> 6.10fF
C6435 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<26> 0.80fF
C6436 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<27> 0.83fF
C6437 BU_3VX2_6|Q BU_3VX2_5|Q 78.85fF
C6438 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<14> 18.82fF
C6439 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<1> 0.44fF
C6440 BU_3VX2_16|Q BU_3VX2_69|Q 1.80fF
C6441 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<15> 21.47fF
C6442 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<13> 12.25fF
C6443 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<8> 3.91fF
C6444 raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<13> 1.64fF
C6445 BU_3VX2_35|Q BU_3VX2_12|Q 1.73fF
C6446 BU_3VX2_64|Q BU_3VX2_9|Q 10.86fF
C6447 BU_3VX2_65|Q BU_3VX2_18|Q 1.91fF
C6448 BU_3VX2_68|Q BU_3VX2_22|Q 14.43fF
C6449 BU_3VX2_69|Q BU_3VX2_30|Q 2.71fF
C6450 BU_3VX2_5|Q BU_3VX2_7|Q 24.36fF
C6451 raven_padframe_0|CORNERESDF_3|VDDR raven_padframe_0|CORNERESDF_3|GNDR 0.68fF
C6452 BU_3VX2_20|A BU_3VX2_17|A 7.28fF
C6453 raven_padframe_0|BBCUD4F_7|VDDR LOGIC0_3V_4|Q 0.01fF
C6454 BU_3VX2_38|A LOGIC0_3V_2|Q 0.03fF
C6455 BU_3VX2_16|A BU_3VX2_27|A 1.90fF
C6456 BU_3VX2_28|A BU_3VX2_14|A 0.01fF
C6457 BU_3VX2_29|A BU_3VX2_27|A 36.13fF
C6458 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<9> 0.01fF
C6459 BU_3VX2_12|A raven_soc_0|flash_csb 0.01fF
C6460 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<10> 23.37fF
C6461 BU_3VX2_73|Q BU_3VX2_46|Q 7.20fF
C6462 raven_soc_0|ram_addr<8> vdd 0.16fF
C6463 raven_soc_0|ram_wdata<22> vdd 0.84fF
C6464 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<11> 0.13fF
C6465 vdd raven_padframe_0|VDDPADF_1|GNDO 0.07fF
C6466 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<11> 0.23fF
C6467 BU_3VX2_37|A BU_3VX2_27|A 0.01fF
C6468 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<14> 0.01fF
C6469 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<9> 1.45fF
C6470 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<13> 0.81fF
C6471 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<7> 0.01fF
C6472 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<6> 0.01fF
C6473 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<12> 22.53fF
C6474 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<27> 12.23fF
C6475 raven_soc_0|ram_rdata<18> raven_soc_0|ram_addr<0> 0.23fF
C6476 raven_soc_0|flash_io1_di raven_soc_0|flash_io2_di 366.95fF
C6477 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<1> 2.56fF
C6478 raven_soc_0|flash_io0_oeb raven_soc_0|flash_io3_di 21.38fF
C6479 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<13> 2.47fF
C6480 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<19> 0.08fF
C6481 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<15> 3.04fF
C6482 BU_3VX2_21|Q BU_3VX2_36|Q 1.40fF
C6483 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<16> 3.69fF
C6484 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io0_di 17.09fF
C6485 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<22> 1.76fF
C6486 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<17> 10.64fF
C6487 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io1_oeb 347.93fF
C6488 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<24> 0.01fF
C6489 raven_soc_0|flash_io1_do raven_soc_0|flash_clk 38.58fF
C6490 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<31> 0.01fF
C6491 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<29> 0.01fF
C6492 raven_soc_0|ram_addr<9> raven_soc_0|ram_addr<2> 4.99fF
C6493 BU_3VX2_36|Q BU_3VX2_8|Q 2.60fF
C6494 LS_3VX2_15|A BU_3VX2_61|Q 169.84fF
C6495 raven_padframe_0|FILLER20F_2|VDDR raven_padframe_0|FILLER20F_2|GNDR 0.68fF
C6496 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<7> 0.01fF
C6497 BU_3VX2_2|A raven_soc_0|flash_io0_di 0.02fF
C6498 BU_3VX2_6|A raven_soc_0|flash_io1_oeb 0.01fF
C6499 raven_soc_0|gpio_pullup<2> raven_soc_0|ext_clk 0.01fF
C6500 BU_3VX2_9|A raven_soc_0|flash_io1_do 0.01fF
C6501 LS_3VX2_11|A LS_3VX2_22|A 12.88fF
C6502 BU_3VX2_38|A raven_soc_0|flash_io0_do 0.01fF
C6503 AMUX4_3V_4|AOUT AMUX4_3V_3|SEL[0] 0.45fF
C6504 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<13> 0.23fF
C6505 LS_3VX2_8|A BU_3VX2_55|Q 0.02fF
C6506 LS_3VX2_5|A BU_3VX2_62|Q 0.01fF
C6507 IN_3VX2_1|A AMUX4_3V_0|SEL[0] 23.24fF
C6508 VDD raven_padframe_0|aregc01_3v3_0|GNDR 0.10fF
C6509 VDD raven_padframe_0|CORNERESDF_0|VDDR 0.71fF
C6510 raven_soc_0|gpio_pulldown<13> BU_3VX2_27|Q 0.01fF
C6511 raven_soc_0|gpio_pulldown<9> apllc03_1v8_0|CLK 0.01fF
C6512 raven_soc_0|gpio_pullup<10> vdd 0.22fF
C6513 raven_soc_0|gpio_outenb<0> BU_3VX2_23|Q 0.01fF
C6514 BU_3VX2_0|Q BU_3VX2_29|Q 0.02fF
C6515 BU_3VX2_20|A BU_3VX2_12|A 2.05fF
C6516 VDD raven_padframe_0|FILLER10F_1|GNDO 0.07fF
C6517 BU_3VX2_35|A raven_soc_0|flash_io2_do 0.08fF
C6518 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<4> 0.01fF
C6519 BU_3VX2_17|A BU_3VX2_14|Q 0.02fF
C6520 BU_3VX2_63|Q raven_soc_0|flash_io3_oeb 0.01fF
C6521 raven_soc_0|gpio_pulldown<0> BU_3VX2_29|Q 0.01fF
C6522 AMUX2_3V_0|SEL AMUX4_3V_1|SEL[1] 8.93fF
C6523 raven_soc_0|gpio_pullup<1> BU_3VX2_27|Q 0.01fF
C6524 BU_3VX2_40|Q raven_soc_0|gpio_in<14> 0.01fF
C6525 BU_3VX2_53|A BU_3VX2_54|A 12.22fF
C6526 BU_3VX2_52|A BU_3VX2_55|A 2.16fF
C6527 VDD3V3 BU_3VX2_57|A 0.05fF
C6528 raven_soc_0|gpio_in<9> VDD3V3 0.07fF
C6529 raven_soc_0|irq_pin BU_3VX2_56|Q 0.01fF
C6530 VDD3V3 BU_3VX2_42|Q 0.02fF
C6531 BU_3VX2_48|Q BU_3VX2_49|Q 211.09fF
C6532 BU_3VX2_3|A BU_3VX2_18|A 0.01fF
C6533 BU_3VX2_15|A BU_3VX2_18|A 7.81fF
C6534 raven_spi_0|SDI raven_spi_0|sdo_enb 13.24fF
C6535 BU_3VX2_23|A BU_3VX2_26|A 11.37fF
C6536 LS_3VX2_14|A LS_3VX2_6|A 14.97fF
C6537 LS_3VX2_3|Q BU_3VX2_27|A 0.01fF
C6538 IN_3VX2_1|A analog_out 1.75fF
C6539 LS_3VX2_7|A AMUX2_3V_0|SEL 18.20fF
C6540 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<8> 0.03fF
C6541 BU_3VX2_31|A raven_soc_0|gpio_pullup<12> 0.01fF
C6542 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<10> 0.01fF
C6543 markings_0|efabless_logo_0|m1_1500_n3150# markings_0|efabless_logo_0|m1_600_n4050# 0.22fF
C6544 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<5> 0.14fF
C6545 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<14> 0.02fF
C6546 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<19> 0.50fF
C6547 raven_soc_0|flash_io0_oeb raven_soc_0|irq_pin 0.54fF
C6548 raven_soc_0|gpio_pullup<6> BU_3VX2_40|Q 0.05fF
C6549 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pullup<5> 4.24fF
C6550 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<13> 0.02fF
C6551 BU_3VX2_6|Q BU_3VX2_28|Q 4.67fF
C6552 BU_3VX2_12|Q BU_3VX2_23|Q 6.21fF
C6553 BU_3VX2_13|Q BU_3VX2_26|Q 2.77fF
C6554 BU_3VX2_38|Q BU_3VX2_25|Q 0.05fF
C6555 BU_3VX2_16|Q BU_3VX2_29|Q 2.67fF
C6556 BU_3VX2_22|Q BU_3VX2_24|Q 23.66fF
C6557 BU_3VX2_67|Q BU_3VX2_25|Q 2.40fF
C6558 BU_3VX2_30|Q BU_3VX2_29|Q 56.86fF
C6559 BU_3VX2_65|Q BU_3VX2_27|Q 0.76fF
C6560 BU_3VX2_7|Q BU_3VX2_28|Q 0.02fF
C6561 BU_3VX2_23|A BU_3VX2_11|A 1.74fF
C6562 raven_soc_0|gpio_outenb<4> BU_3VX2_63|Q 0.20fF
C6563 BU_3VX2_10|A BU_3VX2_7|Q 0.02fF
C6564 LS_3VX2_24|A BU_3VX2_49|Q 6.97fF
C6565 LS_3VX2_4|A BU_3VX2_55|Q 15.41fF
C6566 raven_soc_0|ram_rdata<13> raven_soc_0|ram_rdata<15> 31.52fF
C6567 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<7> 0.02fF
C6568 LS_3VX2_22|A LS_3VX2_21|A 13.99fF
C6569 BU_3VX2_48|A vdd 0.06fF
C6570 AMUX4_3V_1|SEL[1] BU_3VX2_61|Q 8.71fF
C6571 raven_soc_0|flash_io1_oeb BU_3VX2_25|Q 0.01fF
C6572 raven_soc_0|flash_io0_di apllc03_1v8_0|CLK 85.14fF
C6573 raven_soc_0|flash_io0_do BU_3VX2_23|Q 0.01fF
C6574 raven_soc_0|flash_io3_di BU_3VX2_29|Q 0.01fF
C6575 raven_soc_0|flash_io2_di BU_3VX2_28|Q 0.01fF
C6576 raven_padframe_0|FILLER50F_0|VDDR raven_padframe_0|FILLER50F_0|GNDO 0.13fF
C6577 raven_padframe_0|aregc01_3v3_1|VDDR raven_padframe_0|aregc01_3v3_1|GNDO 0.10fF
C6578 raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# raven_padframe_0|axtoc02_3v3_0|GNDR 0.15fF
C6579 markings_0|manufacturer_0|_alphabet_S_1|m2_32_224# markings_0|product_name_0|_alphabet_1_0|m2_64_1376# 0.27fF
C6580 markings_0|mask_copyright_0|m2_n208_960# markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# 0.12fF
C6581 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<12> 0.26fF
C6582 BU_3VX2_10|A raven_soc_0|flash_io2_di 0.04fF
C6583 raven_spi_0|SDI raven_soc_0|gpio_in<15> 2.31fF
C6584 BU_3VX2_63|A raven_soc_0|flash_io0_oeb 0.01fF
C6585 IN_3VX2_1|A raven_soc_0|gpio_in<8> 0.01fF
C6586 BU_3VX2_28|A raven_soc_0|flash_io1_do 4.12fF
C6587 LS_3VX2_7|A BU_3VX2_61|Q 0.01fF
C6588 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<9> 0.07fF
C6589 raven_soc_0|gpio_outenb<15> BU_3VX2_40|Q 2.65fF
C6590 LS_3VX2_6|A BU_3VX2_56|Q 8.63fF
C6591 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<15> 0.02fF
C6592 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<6> 0.01fF
C6593 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pullup<5> 0.02fF
C6594 BU_3VX2_0|Q raven_soc_0|flash_io2_do 0.01fF
C6595 raven_soc_0|gpio_outenb<14> raven_soc_0|ext_clk 0.01fF
C6596 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<14> 0.02fF
C6597 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<11> 28.66fF
C6598 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<19> 0.42fF
C6599 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<23> 12.43fF
C6600 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<20> 8.48fF
C6601 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<28> 0.01fF
C6602 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<0> 1.13fF
C6603 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<15> 0.01fF
C6604 raven_spi_0|CSB raven_soc_0|gpio_out<15> 2.75fF
C6605 BU_3VX2_5|A raven_soc_0|flash_io3_oeb 0.01fF
C6606 BU_3VX2_0|A raven_soc_0|flash_io2_di 12.22fF
C6607 IN_3VX2_1|Q BU_3VX2_59|Q 0.01fF
C6608 IN_3VX2_1|A raven_soc_0|gpio_pullup<13> 0.01fF
C6609 LS_3VX2_10|Q LS_3VX2_19|A 0.01fF
C6610 LS_3VX2_11|A BU_3VX2_60|Q 0.01fF
C6611 VDD raven_padframe_0|BT4F_0|GNDO 0.07fF
C6612 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<9> 7.63fF
C6613 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<8> 0.03fF
C6614 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<14> 0.60fF
C6615 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<27> 0.10fF
C6616 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<29> 0.12fF
C6617 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pullup<6> 16.09fF
C6618 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<10> 0.01fF
C6619 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pulldown<6> 0.02fF
C6620 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<8> 6.65fF
C6621 BU_3VX2_27|A raven_soc_0|flash_io1_oeb 5.79fF
C6622 BU_3VX2_63|Q apllc03_1v8_0|CLK 72.48fF
C6623 raven_soc_0|gpio_pulldown<14> BU_3VX2_23|Q 0.01fF
C6624 raven_soc_0|gpio_pulldown<11> BU_3VX2_28|Q 0.01fF
C6625 raven_padframe_0|BBCUD4F_2|VDDR raven_padframe_0|BBCUD4F_2|VDDO 0.06fF
C6626 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<12> 17.39fF
C6627 BU_3VX2_35|Q BU_3VX2_5|Q 4.63fF
C6628 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<1> 1.82fF
C6629 BU_3VX2_68|Q BU_3VX2_31|Q 0.74fF
C6630 VDD raven_padframe_0|FILLER02F_1|VDDR 0.71fF
C6631 BU_3VX2_2|A BU_3VX2_5|A 3.30fF
C6632 raven_padframe_0|CORNERESDF_2|VDDR raven_padframe_0|CORNERESDF_2|GNDO 0.13fF
C6633 IN_3VX2_1|A BU_3VX2_26|A 8.65fF
C6634 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<14> 0.01fF
C6635 raven_padframe_0|APR00DF_3|GNDR raven_padframe_0|APR00DF_3|GNDO 0.81fF
C6636 raven_padframe_0|FILLER02F_1|VDDO raven_padframe_0|FILLER02F_1|GNDO 2.32fF
C6637 raven_padframe_0|FILLER02F_0|GNDR raven_padframe_0|FILLER02F_0|GNDO 0.84fF
C6638 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<12> 27.89fF
C6639 LS_3VX2_18|A VDD3V3 0.88fF
C6640 raven_soc_0|ram_rdata<27> vdd 0.31fF
C6641 raven_soc_0|ram_wdata<16> apllc03_1v8_0|CLK 0.01fF
C6642 BU_3VX2_3|A BU_3VX2_71|A 0.01fF
C6643 BU_3VX2_15|A BU_3VX2_71|A 0.01fF
C6644 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<11> 0.01fF
C6645 LS_3VX2_10|Q adc_low 0.12fF
C6646 IN_3VX2_1|A BU_3VX2_11|A 0.01fF
C6647 BU_3VX2_65|A BU_3VX2_69|A 3.33fF
C6648 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<8> 1.68fF
C6649 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<2> 1.03fF
C6650 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<4> 0.13fF
C6651 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<15> 0.01fF
C6652 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<12> 158.85fF
C6653 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<15> 0.77fF
C6654 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<12> 38.98fF
C6655 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<14> 1.64fF
C6656 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<9> 0.07fF
C6657 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<11> 0.02fF
C6658 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<6> 0.01fF
C6659 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<13> 0.02fF
C6660 BU_3VX2_7|A raven_soc_0|ext_clk 0.01fF
C6661 raven_soc_0|gpio_pullup<0> VDD3V3 1.46fF
C6662 adc_high VDD3V3 1.54fF
C6663 raven_padframe_0|BBCUD4F_7|VDDR raven_padframe_0|BBCUD4F_7|VDDO 0.06fF
C6664 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<2> 11.63fF
C6665 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<10> 3.24fF
C6666 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<3> 31.18fF
C6667 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<31> 4.40fF
C6668 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<6> 0.01fF
C6669 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<24> 0.01fF
C6670 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<18> 0.01fF
C6671 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<20> 0.01fF
C6672 BU_3VX2_12|Q BU_3VX2_4|Q 4.56fF
C6673 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<26> 15.47fF
C6674 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<29> 0.13fF
C6675 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<1> 0.72fF
C6676 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<25> 57.86fF
C6677 BU_3VX2_19|Q BU_3VX2_36|Q 12.58fF
C6678 BU_3VX2_66|Q BU_3VX2_32|Q 0.85fF
C6679 raven_soc_0|flash_io2_do raven_soc_0|flash_io3_di 123.91fF
C6680 BU_3VX2_13|Q BU_3VX2_11|Q 23.94fF
C6681 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<31> 0.01fF
C6682 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<14> 0.01fF
C6683 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<19> 0.01fF
C6684 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<13> 5.01fF
C6685 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<2> 0.01fF
C6686 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<17> 0.01fF
C6687 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<27> 0.01fF
C6688 BU_3VX2_32|Q BU_3VX2_20|Q 2.65fF
C6689 BU_3VX2_36|Q BU_3VX2_18|Q 3.75fF
C6690 AMUX4_3V_4|SEL[0] BU_3VX2_7|Q 0.01fF
C6691 raven_padframe_0|BBCUD4F_12|VDDO raven_padframe_0|BBCUD4F_12|GNDO 2.28fF
C6692 raven_soc_0|gpio_out<1> BU_3VX2_0|Q 0.01fF
C6693 raven_spi_0|SDO raven_soc_0|flash_io0_oeb 0.37fF
C6694 BU_3VX2_23|A VDD3V3 0.72fF
C6695 BU_3VX2_38|A raven_soc_0|flash_io1_di 0.01fF
C6696 VDD raven_padframe_0|BT4F_2|GNDO 0.07fF
C6697 raven_padframe_0|FILLER50F_2|VDDR raven_padframe_0|FILLER50F_2|GNDO 0.13fF
C6698 LS_3VX2_8|A BU_3VX2_57|Q 0.02fF
C6699 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<7> 0.01fF
C6700 raven_soc_0|gpio_pulldown<13> BU_3VX2_25|Q 0.01fF
C6701 raven_soc_0|gpio_pulldown<4> vdd 0.34fF
C6702 raven_soc_0|gpio_pulldown<10> BU_3VX2_23|Q 0.01fF
C6703 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<0> 45.73fF
C6704 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<10> 0.01fF
C6705 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<6> 1.32fF
C6706 BU_3VX2_14|A raven_soc_0|flash_io1_do 0.01fF
C6707 BU_3VX2_0|Q raven_soc_0|ram_wdata<24> 0.02fF
C6708 raven_soc_0|gpio_out<2> apllc03_1v8_0|CLK 0.01fF
C6709 raven_soc_0|gpio_pullup<1> BU_3VX2_25|Q 0.01fF
C6710 BU_3VX2_43|A LS_3VX2_20|Q 2.83fF
C6711 BU_3VX2_44|A LS_3VX2_21|Q 0.45fF
C6712 raven_padframe_0|BT4F_1|VDDO raven_padframe_0|BT4F_1|GNDO 2.28fF
C6713 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<6> 0.27fF
C6714 BU_3VX2_31|A raven_soc_0|gpio_outenb<0> 0.01fF
C6715 BU_3VX2_37|A BU_3VX2_37|Q 0.08fF
C6716 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<4> 0.29fF
C6717 raven_padframe_0|BBCUD4F_1|VDDO raven_padframe_0|BBCUD4F_1|GNDO 2.28fF
C6718 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<10> 0.24fF
C6719 LOGIC0_3V_4|Q raven_padframe_0|BBC4F_2|PO 0.04fF
C6720 raven_soc_0|flash_csb raven_soc_0|flash_clk 418.79fF
C6721 BU_3VX2_63|Q raven_soc_0|gpio_outenb<8> 0.01fF
C6722 raven_padframe_0|FILLER10F_0|VDDR raven_padframe_0|FILLER10F_0|VDDO 0.06fF
C6723 BU_3VX2_6|Q vdd 1.35fF
C6724 BU_3VX2_35|Q BU_3VX2_28|Q 0.01fF
C6725 BU_3VX2_7|Q vdd 1.02fF
C6726 BU_3VX2_55|Q vdd 1.77fF
C6727 BU_3VX2_5|Q BU_3VX2_23|Q 8.08fF
C6728 BU_3VX2_65|Q BU_3VX2_25|Q 0.09fF
C6729 BU_3VX2_69|Q BU_3VX2_26|Q 0.01fF
C6730 BU_3VX2_31|Q BU_3VX2_24|Q 4.07fF
C6731 BU_3VX2_68|Q apllc03_1v8_0|CLK 0.91fF
C6732 BU_3VX2_25|A BU_3VX2_26|A 56.38fF
C6733 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<10> 0.01fF
C6734 BU_3VX2_9|A raven_soc_0|flash_csb 0.01fF
C6735 BU_3VX2_68|A VDD3V3 0.02fF
C6736 BU_3VX2_70|A BU_3VX2_68|Q 0.03fF
C6737 LS_3VX2_4|A BU_3VX2_57|Q 11.78fF
C6738 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pulldown<3> 1.53fF
C6739 raven_soc_0|ram_wdata<27> raven_soc_0|ram_rdata<17> 1.08fF
C6740 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<16> 0.01fF
C6741 raven_soc_0|flash_io2_di vdd 5.08fF
C6742 BU_3VX2_1|Q BU_3VX2_52|Q 0.44fF
C6743 BU_3VX2_59|A BU_3VX2_59|Q 0.10fF
C6744 AMUX4_3V_1|SEL[1] LS_3VX2_15|A 8.10fF
C6745 raven_soc_0|flash_io3_oeb BU_3VX2_24|Q 0.01fF
C6746 LS_3VX2_22|A LS_3VX2_27|A 18.36fF
C6747 raven_soc_0|flash_io1_di BU_3VX2_23|Q 0.01fF
C6748 raven_soc_0|flash_io0_oeb BU_3VX2_26|Q 0.01fF
C6749 AMUX4_3V_0|AOUT vdd 0.94fF
C6750 BU_3VX2_49|A BU_3VX2_50|Q 0.03fF
C6751 raven_padframe_0|BT4FC_0|GNDR raven_padframe_0|BT4FC_0|VDDO 0.09fF
C6752 raven_padframe_0|FILLER01F_0|GNDR raven_padframe_0|FILLER01F_0|VDDO 0.09fF
C6753 BU_3VX2_25|A BU_3VX2_11|A 0.01fF
C6754 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<8> 0.01fF
C6755 LOGIC0_3V_4|Q raven_soc_0|gpio_in<4> 0.08fF
C6756 raven_padframe_0|aregc01_3v3_1|m4_92500_22024# raven_padframe_0|aregc01_3v3_1|VDDO 1.17fF
C6757 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<3> 14.32fF
C6758 raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# raven_padframe_0|axtoc02_3v3_0|m4_55000_22024# 0.02fF
C6759 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<9> 0.35fF
C6760 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<12> 0.02fF
C6761 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<11> 0.01fF
C6762 BU_3VX2_8|A BU_3VX2_9|Q 0.03fF
C6763 BU_3VX2_63|A raven_soc_0|flash_io2_do 0.01fF
C6764 BU_3VX2_66|A BU_3VX2_67|Q 0.03fF
C6765 BU_3VX2_18|A BU_3VX2_17|Q 0.16fF
C6766 IN_3VX2_1|A VDD3V3 7.65fF
C6767 LS_3VX2_7|A LS_3VX2_15|A 0.31fF
C6768 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<5> 0.42fF
C6769 LS_3VX2_3|A raven_soc_0|flash_io1_do 0.06fF
C6770 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<15> 0.02fF
C6771 raven_soc_0|gpio_pullup<15> raven_soc_0|ext_clk 0.01fF
C6772 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<14> 0.02fF
C6773 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<12> 0.02fF
C6774 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<9> 17.97fF
C6775 VDD raven_padframe_0|APR00DF_0|GNDR 0.16fF
C6776 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<23> 4.41fF
C6777 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<0> 0.57fF
C6778 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<19> 0.01fF
C6779 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<20> 8.49fF
C6780 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<11> 3.25fF
C6781 BU_3VX2_71|Q BU_3VX2_27|Q 2.44fF
C6782 BU_3VX2_36|Q BU_3VX2_27|Q 8.38fF
C6783 BU_3VX2_10|A BU_3VX2_38|A 0.66fF
C6784 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<7> 0.01fF
C6785 BU_3VX2_20|A raven_soc_0|flash_clk 1.60fF
C6786 LS_3VX2_11|A BU_3VX2_62|Q 0.01fF
C6787 IN_3VX2_1|Q BU_3VX2_61|Q 0.01fF
C6788 LS_3VX2_10|Q LS_3VX2_22|A 0.01fF
C6789 BU_3VX2_40|A raven_soc_0|flash_io2_di 0.48fF
C6790 LOGIC0_3V_4|Q raven_soc_0|gpio_in<7> 0.08fF
C6791 raven_soc_0|gpio_in<2> raven_soc_0|flash_io2_di 0.23fF
C6792 raven_spi_0|sdo_enb raven_soc_0|flash_io0_di 7.39fF
C6793 BU_3VX2_31|A raven_soc_0|flash_io0_do 6.92fF
C6794 BU_3VX2_13|A raven_soc_0|flash_io3_oeb 0.01fF
C6795 LS_3VX2_8|A LS_3VX2_16|A 0.01fF
C6796 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<6> 1.01fF
C6797 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_out<8> 0.08fF
C6798 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<13> 0.01fF
C6799 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<15> 0.01fF
C6800 BU_3VX2_0|Q BU_3VX2_32|Q 0.01fF
C6801 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pulldown<6> 0.02fF
C6802 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<13> 0.02fF
C6803 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pulldown<7> 0.33fF
C6804 VDD raven_padframe_0|axtoc02_3v3_0|VDDR 1.07fF
C6805 raven_soc_0|gpio_pulldown<11> vdd 0.15fF
C6806 LS_3VX2_13|A BU_3VX2_51|Q 5.56fF
C6807 BU_3VX2_32|A LS_3VX2_2|Q 0.01fF
C6808 BU_3VX2_9|A BU_3VX2_20|A 1.11fF
C6809 BU_3VX2_38|A BU_3VX2_0|A 0.01fF
C6810 BU_3VX2_2|A BU_3VX2_13|A 1.32fF
C6811 LS_3VX2_11|A LS_3VX2_5|A 34.88fF
C6812 raven_padframe_0|ICFC_0|VDDR raven_padframe_0|ICFC_0|GNDO 0.13fF
C6813 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<8> 0.44fF
C6814 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_out<14> 0.18fF
C6815 BU_3VX2_24|A BU_3VX2_3|A 0.01fF
C6816 BU_3VX2_24|A BU_3VX2_15|A 2.29fF
C6817 BU_3VX2_53|A BU_3VX2_53|Q 0.10fF
C6818 LS_3VX2_12|A LS_3VX2_10|A 23.14fF
C6819 LS_3VX2_13|Q LS_3VX2_11|Q 2.01fF
C6820 raven_spi_0|SDI raven_soc_0|gpio_outenb<15> 2.95fF
C6821 BU_3VX2_31|A raven_soc_0|gpio_pulldown<14> 0.01fF
C6822 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<11> 0.01fF
C6823 BU_3VX2_28|A raven_soc_0|flash_csb 12.74fF
C6824 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<11> 11.15fF
C6825 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<14> 0.09fF
C6826 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<12> 58.85fF
C6827 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<10> 0.04fF
C6828 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<15> 0.02fF
C6829 BU_3VX2_0|Q raven_soc_0|gpio_out<11> 0.01fF
C6830 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<13> 0.02fF
C6831 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<18> 6.78fF
C6832 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<24> 34.58fF
C6833 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<30> 2.02fF
C6834 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<23> 0.26fF
C6835 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<6> 6.62fF
C6836 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<31> 0.14fF
C6837 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<20> 10.62fF
C6838 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<21> 4.47fF
C6839 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<9> 0.02fF
C6840 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<22> 0.01fF
C6841 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<7> 3.95fF
C6842 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<3> 0.01fF
C6843 BU_3VX2_38|Q BU_3VX2_37|Q 65.59fF
C6844 BU_3VX2_4|Q BU_3VX2_5|Q 74.77fF
C6845 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<8> 0.05fF
C6846 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<12> 26.12fF
C6847 BU_3VX2_70|Q BU_3VX2_7|Q 0.40fF
C6848 BU_3VX2_12|Q BU_3VX2_3|Q 9.33fF
C6849 BU_3VX2_14|Q BU_3VX2_10|Q 9.86fF
C6850 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<21> 0.11fF
C6851 BU_3VX2_2|Q BU_3VX2_14|Q 2.75fF
C6852 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<17> 0.02fF
C6853 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<2> 12.74fF
C6854 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<2> 6.39fF
C6855 BU_3VX2_6|Q BU_3VX2_70|Q 2.56fF
C6856 BU_3VX2_11|Q BU_3VX2_69|Q 0.01fF
C6857 BU_3VX2_32|Q BU_3VX2_30|Q 1.07fF
C6858 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<13> 5.07fF
C6859 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<25> 5.97fF
C6860 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<26> 0.03fF
C6861 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<19> 4.93fF
C6862 BU_3VX2_43|Q BU_3VX2_46|Q 49.76fF
C6863 BU_3VX2_42|Q adc0_data<5> 19.21fF
C6864 BU_3VX2_23|Q BU_3VX2_28|Q 56.11fF
C6865 BU_3VX2_26|Q BU_3VX2_29|Q 91.03fF
C6866 BU_3VX2_24|Q apllc03_1v8_0|CLK 1.05fF
C6867 raven_padframe_0|FILLER50F_1|VDDR raven_padframe_0|FILLER50F_1|GNDR 0.68fF
C6868 raven_padframe_0|CORNERESDF_0|GNDR raven_padframe_0|CORNERESDF_0|GNDO 0.81fF
C6869 LOGIC0_3V_4|Q raven_soc_0|gpio_out<7> 0.01fF
C6870 raven_spi_0|SDO raven_soc_0|flash_io2_do 0.62fF
C6871 raven_padframe_0|FILLER20F_1|VDDR raven_padframe_0|FILLER20F_1|VDDO 0.06fF
C6872 LS_3VX2_7|A AMUX4_3V_1|SEL[1] 12.25fF
C6873 LS_3VX2_4|A LS_3VX2_16|A 0.09fF
C6874 BU_3VX2_64|A BU_3VX2_65|Q 0.03fF
C6875 raven_soc_0|gpio_pulldown<12> BU_3VX2_23|Q 0.01fF
C6876 BU_3VX2_71|Q raven_soc_0|flash_io2_oeb 0.05fF
C6877 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<13> 9.27fF
C6878 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<15> 11.69fF
C6879 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<17> 0.37fF
C6880 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<1> 0.10fF
C6881 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<16> 5.42fF
C6882 raven_soc_0|ram_rdata<20> raven_soc_0|ram_addr<0> 4.30fF
C6883 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<12> 0.01fF
C6884 BU_3VX2_37|A BU_3VX2_40|Q 0.02fF
C6885 BU_3VX2_25|A VDD3V3 0.54fF
C6886 raven_soc_0|gpio_out<3> raven_soc_0|ext_clk 0.01fF
C6887 VDD raven_padframe_0|aregc01_3v3_1|GNDO 0.06fF
C6888 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<11> 148.18fF
C6889 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<12> 0.01fF
C6890 BU_3VX2_63|Q raven_soc_0|gpio_in<15> 0.01fF
C6891 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<5> 0.01fF
C6892 BU_3VX2_20|A BU_3VX2_28|A 2.66fF
C6893 BU_3VX2_4|A BU_3VX2_26|A 0.01fF
C6894 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<8> 0.11fF
C6895 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<4> 0.02fF
C6896 BU_3VX2_22|A raven_soc_0|flash_io0_do 0.01fF
C6897 BU_3VX2_31|A raven_soc_0|gpio_pulldown<10> 0.01fF
C6898 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_outenb<0> 4.27fF
C6899 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<8> 0.01fF
C6900 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<9> 4.94fF
C6901 BU_3VX2_35|Q vdd 0.35fF
C6902 BU_3VX2_57|Q vdd 1.89fF
C6903 LS_3VX2_23|Q BU_3VX2_32|A 8.23fF
C6904 VDD3V3 raven_padframe_0|VDDPADFC_0|GNDR 0.16fF
C6905 BU_3VX2_3|A BU_3VX2_16|A 0.75fF
C6906 BU_3VX2_16|A BU_3VX2_15|A 39.08fF
C6907 BU_3VX2_3|A BU_3VX2_29|A 0.01fF
C6908 LS_3VX2_5|Q LS_3VX2_9|Q 8.07fF
C6909 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<4> 0.64fF
C6910 BU_3VX2_4|A BU_3VX2_11|A 1.49fF
C6911 BU_3VX2_15|A BU_3VX2_29|A 0.01fF
C6912 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_outenb<2> 22.73fF
C6913 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<13> 0.01fF
C6914 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<17> 0.02fF
C6915 LS_3VX2_22|A BU_3VX2_1|Q 0.10fF
C6916 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<27> 0.01fF
C6917 raven_soc_0|ram_wdata<22> raven_soc_0|ram_wdata<27> 21.47fF
C6918 raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<15> 2.09fF
C6919 raven_soc_0|ram_wdata<25> raven_soc_0|ram_wdata<31> 17.18fF
C6920 raven_soc_0|ram_wdata<21> raven_soc_0|ram_rdata<1> 1.45fF
C6921 raven_soc_0|ram_wdata<26> raven_soc_0|ram_rdata<17> 0.02fF
C6922 raven_soc_0|ram_wdata<17> raven_soc_0|ram_addr<0> 0.01fF
C6923 BU_3VX2_49|A LS_3VX2_27|Q 0.11fF
C6924 BU_3VX2_48|A LS_3VX2_21|Q 0.15fF
C6925 BU_3VX2_47|A BU_3VX2_43|A 0.47fF
C6926 raven_soc_0|gpio_out<15> apllc03_1v8_0|CLK 0.01fF
C6927 BU_3VX2_59|A BU_3VX2_61|Q 0.03fF
C6928 LS_3VX2_17|Q BU_3VX2_62|Q 0.23fF
C6929 LS_3VX2_19|A BU_3VX2_53|Q 6.56fF
C6930 raven_soc_0|flash_io2_do BU_3VX2_26|Q 0.01fF
C6931 BU_3VX2_53|Q BU_3VX2_52|Q 228.31fF
C6932 BU_3VX2_46|Q BU_3VX2_50|Q 27.76fF
C6933 BU_3VX2_49|A BU_3VX2_48|Q 0.15fF
C6934 BU_3VX2_3|A BU_3VX2_37|A 5.40fF
C6935 raven_padframe_0|aregc01_3v3_1|m4_0_29057# raven_padframe_0|aregc01_3v3_1|VDDO 0.04fF
C6936 raven_padframe_0|aregc01_3v3_1|m4_0_29333# raven_padframe_0|aregc01_3v3_1|GNDO 0.12fF
C6937 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<1> 0.17fF
C6938 raven_padframe_0|axtoc02_3v3_0|m4_55000_30653# raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# 0.03fF
C6939 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<12> 0.02fF
C6940 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<6> 0.01fF
C6941 BU_3VX2_14|A raven_soc_0|flash_csb 0.01fF
C6942 BU_3VX2_63|Q raven_soc_0|gpio_out<13> 0.01fF
C6943 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<10> 0.01fF
C6944 markings_0|date_0|_alphabet_1_1|m2_64_1376# markings_0|date_0|_alphabet_2_0|m2_0_0# 0.03fF
C6945 markings_0|mask_copyright_0|m2_n208_960# markings_0|mask_copyright_0|m2_1056_1056# 0.77fF
C6946 BU_3VX2_38|A vdd 0.27fF
C6947 BU_3VX2_40|A BU_3VX2_35|Q 0.03fF
C6948 BU_3VX2_66|A BU_3VX2_65|Q 0.16fF
C6949 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<7> 0.01fF
C6950 BU_3VX2_0|Q raven_soc_0|gpio_in<12> 0.01fF
C6951 LS_3VX2_3|A raven_soc_0|gpio_in<10> 0.17fF
C6952 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<8> 0.02fF
C6953 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<14> 0.02fF
C6954 raven_soc_0|gpio_pullup<3> VDD3V3 0.23fF
C6955 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<28> 16.99fF
C6956 raven_padframe_0|FILLER02F_1|VDDR raven_padframe_0|FILLER02F_1|GNDR 0.68fF
C6957 BU_3VX2_4|Q BU_3VX2_28|Q 2.63fF
C6958 BU_3VX2_36|Q BU_3VX2_25|Q 1.97fF
C6959 BU_3VX2_11|Q BU_3VX2_29|Q 0.01fF
C6960 raven_soc_0|gpio_pullup<14> BU_3VX2_27|Q 0.01fF
C6961 raven_soc_0|gpio_outenb<13> BU_3VX2_29|Q 0.01fF
C6962 BU_3VX2_71|Q BU_3VX2_25|Q 2.02fF
C6963 raven_soc_0|gpio_in<5> apllc03_1v8_0|CLK 0.01fF
C6964 LS_3VX2_23|A apllc03_1v8_0|CLK 2.01fF
C6965 LS_3VX2_21|A BU_3VX2_45|Q 8.81fF
C6966 BU_3VX2_23|A BU_3VX2_21|Q 0.03fF
C6967 AMUX4_3V_0|AIN1 BU_3VX2_42|Q 0.14fF
C6968 IN_3VX2_1|Q LS_3VX2_15|A 0.01fF
C6969 aporc02_3v3_0|PORB VDD3V3 0.10fF
C6970 VDD raven_padframe_0|VDDORPADF_4|GNDO 0.07fF
C6971 BU_3VX2_18|A raven_soc_0|flash_io0_di 0.01fF
C6972 raven_padframe_0|BBC4F_3|VDDR raven_padframe_0|BBC4F_3|VDDO 0.06fF
C6973 BU_3VX2_31|A raven_soc_0|flash_io1_di 3.70fF
C6974 VDD raven_padframe_0|FILLER50F_0|VDDR 0.71fF
C6975 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<1> 15.82fF
C6976 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pulldown<7> 75.12fF
C6977 VDD raven_padframe_0|BBCUD4F_9|GNDO 0.07fF
C6978 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<15> 0.26fF
C6979 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<9> 4.31fF
C6980 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<0> 9.18fF
C6981 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pulldown<3> 0.68fF
C6982 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<5> 19.14fF
C6983 BU_3VX2_33|A raven_soc_0|flash_io3_do 0.21fF
C6984 adc_low BU_3VX2_53|Q 0.05fF
C6985 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pulldown<6> 0.01fF
C6986 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<13> 0.02fF
C6987 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<6> 0.01fF
C6988 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<8> 3.20fF
C6989 BU_3VX2_0|Q raven_soc_0|ram_rdata<16> 0.02fF
C6990 LS_3VX2_13|A BU_3VX2_49|Q 4.69fF
C6991 raven_padframe_0|FILLER02F_0|VDDR raven_padframe_0|FILLER02F_0|GNDO 0.13fF
C6992 BU_3VX2_46|A BU_3VX2_45|A 6.92fF
C6993 BU_3VX2_38|A BU_3VX2_40|A 8.89fF
C6994 BU_3VX2_21|A raven_soc_0|flash_io0_do 0.01fF
C6995 LS_3VX2_12|A raven_soc_0|ser_tx 0.01fF
C6996 BU_3VX2_38|Q BU_3VX2_40|Q 0.21fF
C6997 BU_3VX2_55|A BU_3VX2_55|Q 0.10fF
C6998 raven_soc_0|irq_pin AMUX4_3V_4|AIN2 12.56fF
C6999 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<4> 0.01fF
C7000 BU_3VX2_23|A BU_3VX2_19|A 5.63fF
C7001 BU_3VX2_3|A LS_3VX2_3|Q 0.01fF
C7002 LS_3VX2_12|A LS_3VX2_24|A 14.93fF
C7003 LS_3VX2_3|Q BU_3VX2_15|A 0.01fF
C7004 AMUX4_3V_4|AOUT AMUX4_3V_4|AIN1 0.37fF
C7005 BU_3VX2_20|A BU_3VX2_14|A 3.00fF
C7006 IN_3VX2_1|A raven_soc_0|gpio_pullup<8> 0.01fF
C7007 raven_soc_0|gpio_in<0> LS_3VX2_3|A 0.01fF
C7008 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_outenb<5> 0.04fF
C7009 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<12> 28.73fF
C7010 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<15> 0.90fF
C7011 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<11> 0.52fF
C7012 LS_3VX2_3|A raven_soc_0|flash_csb 0.01fF
C7013 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<14> 0.01fF
C7014 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<15> 0.02fF
C7015 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<5> 0.07fF
C7016 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<6> 0.01fF
C7017 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<7> 0.01fF
C7018 raven_soc_0|gpio_out<1> BU_3VX2_26|Q 0.01fF
C7019 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<23> 4.44fF
C7020 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<14> 0.36fF
C7021 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<7> 6.84fF
C7022 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<30> 1.53fF
C7023 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<21> 0.12fF
C7024 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<4> 0.21fF
C7025 BU_3VX2_3|Q BU_3VX2_5|Q 47.01fF
C7026 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<25> 11.59fF
C7027 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<14> 5.14fF
C7028 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<2> 0.01fF
C7029 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<12> 0.01fF
C7030 BU_3VX2_40|Q raven_soc_0|flash_io1_oeb 0.18fF
C7031 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<15> 0.01fF
C7032 LS_3VX2_16|A vdd 1.53fF
C7033 AMUX4_3V_0|SEL[1] BU_3VX2_72|Q 0.77fF
C7034 vdd BU_3VX2_23|Q 0.78fF
C7035 BU_3VX2_51|Q BU_3VX2_72|Q 3.24fF
C7036 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<2> 5.73fF
C7037 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<11> 0.01fF
C7038 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<7> 0.01fF
C7039 raven_padframe_0|aregc01_3v3_0|m4_92500_22024# raven_padframe_0|aregc01_3v3_0|VDDO 1.17fF
C7040 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<13> 0.12fF
C7041 AMUX4_3V_1|AIN1 BU_3VX2_60|A 0.02fF
C7042 BU_3VX2_4|A VDD3V3 0.25fF
C7043 raven_soc_0|gpio_out<4> vdd 0.20fF
C7044 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<19> 0.01fF
C7045 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<20> 0.01fF
C7046 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<23> 0.01fF
C7047 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_out<15> 0.02fF
C7048 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<22> 1.43fF
C7049 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<29> 0.03fF
C7050 BU_3VX2_1|Q BU_3VX2_60|Q 0.12fF
C7051 raven_soc_0|ram_wdata<20> apllc03_1v8_0|CLK 0.01fF
C7052 BU_3VX2_58|Q BU_3VX2_53|Q 26.91fF
C7053 BU_3VX2_3|A BU_3VX2_38|Q 0.02fF
C7054 AMUX4_3V_0|AIN1 BU_3VX2_42|A 0.45fF
C7055 IN_3VX2_1|Q AMUX4_3V_1|SEL[1] 0.01fF
C7056 AMUX4_3V_4|AOUT VDD3V3 5.78fF
C7057 raven_padframe_0|ICFC_0|VDD3 raven_padframe_0|ICFC_0|GNDO 0.07fF
C7058 BU_3VX2_26|A raven_soc_0|flash_io0_oeb 4.06fF
C7059 BU_3VX2_31|A BU_3VX2_28|Q 81.84fF
C7060 BU_3VX2_63|Q raven_soc_0|gpio_in<14> 0.01fF
C7061 raven_soc_0|gpio_in<2> BU_3VX2_23|Q 0.01fF
C7062 BU_3VX2_0|Q raven_soc_0|ram_rdata<22> 0.02fF
C7063 AMUX2_3V_0|SEL LS_3VX2_20|A 8.21fF
C7064 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<10> 0.11fF
C7065 raven_soc_0|gpio_in<5> raven_soc_0|gpio_outenb<8> 0.01fF
C7066 raven_padframe_0|FILLER10F_1|GNDR raven_padframe_0|FILLER10F_1|GNDO 0.81fF
C7067 BU_3VX2_10|A BU_3VX2_31|A 0.01fF
C7068 BU_3VX2_31|A raven_soc_0|gpio_pulldown<12> 0.01fF
C7069 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<2> 1.77fF
C7070 BU_3VX2_22|A raven_soc_0|flash_io1_di 0.01fF
C7071 BU_3VX2_3|A raven_soc_0|flash_io1_oeb 0.01fF
C7072 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<10> 0.01fF
C7073 BU_3VX2_15|A raven_soc_0|flash_io1_oeb 0.01fF
C7074 LS_3VX2_11|Q LS_3VX2_19|A 0.01fF
C7075 BU_3VX2_71|A raven_soc_0|flash_io0_di 0.01fF
C7076 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<10> 0.01fF
C7077 raven_soc_0|gpio_in<3> raven_soc_0|flash_io3_oeb 0.93fF
C7078 BU_3VX2_14|A BU_3VX2_14|Q 0.08fF
C7079 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<6> 0.10fF
C7080 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<7> 3.45fF
C7081 BU_3VX2_63|Q raven_soc_0|gpio_pullup<6> 0.05fF
C7082 BU_3VX2_64|A BU_3VX2_36|Q 0.16fF
C7083 IN_3VX2_1|A adc0_data<5> 7.52fF
C7084 BU_3VX2_11|A raven_soc_0|flash_io0_oeb 0.01fF
C7085 raven_soc_0|flash_csb raven_soc_0|flash_io1_do 23.47fF
C7086 BU_3VX2_19|A IN_3VX2_1|A 1.90fF
C7087 BU_3VX2_5|A BU_3VX2_18|A 0.81fF
C7088 BU_3VX2_0|A BU_3VX2_31|A 0.89fF
C7089 BU_3VX2_35|A BU_3VX2_12|A 1.00fF
C7090 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<8> 11.49fF
C7091 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<27> 0.68fF
C7092 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<31> 0.25fF
C7093 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<1> 11.57fF
C7094 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<15> 0.08fF
C7095 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<25> 0.01fF
C7096 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<26> 0.01fF
C7097 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<17> 0.01fF
C7098 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<22> 0.01fF
C7099 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<21> 0.01fF
C7100 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<17> 0.01fF
C7101 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<0> 0.01fF
C7102 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<25> 15.97fF
C7103 LS_3VX2_2|A BU_3VX2_7|Q 0.04fF
C7104 raven_soc_0|ram_wdata<15> raven_soc_0|ram_rdata<13> 0.24fF
C7105 raven_soc_0|ram_wdata<14> raven_soc_0|ram_rdata<1> 0.33fF
C7106 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<22> 25.30fF
C7107 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<31> 0.01fF
C7108 LS_3VX2_22|A BU_3VX2_53|Q 0.02fF
C7109 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<29> 6.14fF
C7110 raven_soc_0|gpio_in<6> apllc03_1v8_0|CLK 0.02fF
C7111 raven_soc_0|gpio_in<8> BU_3VX2_29|Q 0.01fF
C7112 raven_soc_0|gpio_in<15> BU_3VX2_24|Q 0.01fF
C7113 raven_soc_0|gpio_in<11> BU_3VX2_23|Q 0.01fF
C7114 raven_soc_0|gpio_in<9> BU_3VX2_27|Q 0.01fF
C7115 BU_3VX2_46|Q BU_3VX2_48|Q 46.28fF
C7116 raven_spi_0|SDI BU_3VX2_37|A 0.17fF
C7117 raven_padframe_0|VDDPADFC_0|VDDO raven_padframe_0|VDDPADFC_0|GNDO 2.28fF
C7118 LS_3VX2_11|Q adc_low 0.12fF
C7119 raven_padframe_0|aregc01_3v3_1|m4_92500_29057# raven_padframe_0|aregc01_3v3_1|m4_92500_28769# 0.11fF
C7120 BU_3VX2_71|A BU_3VX2_63|Q 0.03fF
C7121 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_in<3> 2.73fF
C7122 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<10> 0.01fF
C7123 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<11> 0.01fF
C7124 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<14> 7.23fF
C7125 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<12> 0.02fF
C7126 BU_3VX2_63|Q raven_soc_0|gpio_outenb<15> 0.01fF
C7127 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<13> 0.34fF
C7128 BU_3VX2_7|A BU_3VX2_7|Q 0.08fF
C7129 BU_3VX2_7|A BU_3VX2_6|Q 0.16fF
C7130 LS_3VX2_14|A VDD3V3 0.48fF
C7131 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<11> 0.39fF
C7132 raven_soc_0|gpio_pulldown<13> BU_3VX2_40|Q 0.03fF
C7133 LS_3VX2_3|A raven_soc_0|gpio_in<13> 0.95fF
C7134 raven_soc_0|gpio_pulldown<5> VDD3V3 0.30fF
C7135 BU_3VX2_3|Q BU_3VX2_28|Q 0.27fF
C7136 BU_3VX2_4|Q vdd 1.37fF
C7137 BU_3VX2_32|Q BU_3VX2_26|Q 1.58fF
C7138 BU_3VX2_70|Q BU_3VX2_23|Q 5.65fF
C7139 raven_soc_0|gpio_pullup<14> BU_3VX2_25|Q 0.01fF
C7140 raven_soc_0|gpio_pullup<13> BU_3VX2_29|Q 0.01fF
C7141 raven_soc_0|gpio_out<8> BU_3VX2_28|Q 0.01fF
C7142 raven_soc_0|gpio_out<10> apllc03_1v8_0|CLK 0.01fF
C7143 LS_3VX2_27|A BU_3VX2_45|Q 7.95fF
C7144 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<4> 52.70fF
C7145 BU_3VX2_7|A raven_soc_0|flash_io2_di 0.01fF
C7146 BU_3VX2_8|A raven_soc_0|flash_io3_do 0.01fF
C7147 BU_3VX2_20|A raven_soc_0|flash_io1_do 0.01fF
C7148 BU_3VX2_17|A BU_3VX2_16|Q 0.16fF
C7149 BU_3VX2_16|A BU_3VX2_17|Q 0.03fF
C7150 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<9> 0.10fF
C7151 raven_soc_0|gpio_pullup<1> BU_3VX2_40|Q 0.04fF
C7152 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pulldown<6> 0.69fF
C7153 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<14> 0.28fF
C7154 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<5> 0.01fF
C7155 BU_3VX2_0|Q raven_soc_0|gpio_pulldown<7> 0.26fF
C7156 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<8> 0.01fF
C7157 LS_3VX2_24|A BU_3VX2_46|Q 4.78fF
C7158 raven_spi_0|sdo_enb raven_soc_0|gpio_out<15> 1.53fF
C7159 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<23> 18.18fF
C7160 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<19> 5.11fF
C7161 BU_3VX2_49|A BU_3VX2_41|A 1.72fF
C7162 BU_3VX2_50|A BU_3VX2_46|A 0.84fF
C7163 raven_padframe_0|APR00DF_6|GNDR raven_padframe_0|APR00DF_6|GNDO 0.81fF
C7164 BU_3VX2_21|A raven_soc_0|flash_io1_di 0.13fF
C7165 BU_3VX2_17|A raven_soc_0|flash_io3_di 0.01fF
C7166 LS_3VX2_11|A LS_3VX2_21|A 5.36fF
C7167 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<7> 1.34fF
C7168 BU_3VX2_66|A BU_3VX2_36|Q 0.02fF
C7169 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<6> 0.01fF
C7170 raven_soc_0|ram_wdata<3> vdd 1.01fF
C7171 raven_soc_0|gpio_out<9> apllc03_1v8_0|CLK 0.01fF
C7172 raven_soc_0|gpio_in<3> apllc03_1v8_0|CLK 0.01fF
C7173 raven_soc_0|gpio_out<13> BU_3VX2_24|Q 0.01fF
C7174 raven_soc_0|gpio_out<11> BU_3VX2_26|Q 0.01fF
C7175 BU_3VX2_73|Q raven_soc_0|ext_clk 0.01fF
C7176 BU_3VX2_55|A BU_3VX2_57|Q 0.04fF
C7177 BU_3VX2_10|A BU_3VX2_22|A 1.31fF
C7178 LS_3VX2_12|Q LS_3VX2_9|Q 0.74fF
C7179 raven_padframe_0|axtoc02_3v3_0|XI XI 2.38fF
C7180 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<7> 0.01fF
C7181 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<7> 1.10fF
C7182 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<11> 0.52fF
C7183 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<8> 0.38fF
C7184 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<6> 4.40fF
C7185 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<11> 30.37fF
C7186 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<6> 0.01fF
C7187 raven_soc_0|gpio_in<4> BU_3VX2_71|Q 0.02fF
C7188 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<6> 0.01fF
C7189 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<6> 5.37fF
C7190 AMUX2_3V_0|SEL BU_3VX2_47|Q 4.75fF
C7191 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<1> 0.01fF
C7192 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<12> 1.07fF
C7193 raven_soc_0|gpio_in<15> raven_soc_0|gpio_out<15> 117.52fF
C7194 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<7> 0.17fF
C7195 raven_soc_0|ext_clk raven_soc_0|flash_io3_oeb 16.94fF
C7196 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<5> 0.01fF
C7197 raven_soc_0|flash_io0_oeb VDD3V3 12.73fF
C7198 BU_3VX2_49|Q BU_3VX2_72|Q 6.47fF
C7199 VDD raven_padframe_0|FILLER40F_0|VDDR 0.71fF
C7200 BU_3VX2_19|A BU_3VX2_25|A 3.60fF
C7201 BU_3VX2_22|A BU_3VX2_0|A 0.01fF
C7202 raven_spi_0|SDI LOGIC0_3V_4|Q 1.02fF
C7203 BU_3VX2_5|A BU_3VX2_71|A 0.01fF
C7204 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<9> 0.01fF
C7205 raven_padframe_0|aregc01_3v3_0|m4_92500_29333# raven_padframe_0|aregc01_3v3_0|m4_92500_22024# 0.01fF
C7206 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<15> 0.69fF
C7207 AMUX4_3V_1|AIN1 VDD3V3 2.18fF
C7208 BU_3VX2_2|A raven_soc_0|ext_clk 0.02fF
C7209 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<2> 0.22fF
C7210 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<0> 0.96fF
C7211 BU_3VX2_71|Q raven_soc_0|gpio_in<7> 0.45fF
C7212 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<20> 9.40fF
C7213 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<21> 0.01fF
C7214 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<6> 1.65fF
C7215 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<15> 0.01fF
C7216 raven_soc_0|ram_addr<2> vdd 0.22fF
C7217 BU_3VX2_60|Q BU_3VX2_53|Q 18.43fF
C7218 raven_soc_0|ram_rdata<21> apllc03_1v8_0|CLK 0.01fF
C7219 raven_padframe_0|FILLER40F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C7220 AMUX4_3V_3|AOUT AMUX4_3V_3|SEL[0] 0.26fF
C7221 LS_3VX2_9|A BU_3VX2_55|Q 13.47fF
C7222 BU_3VX2_12|A raven_soc_0|flash_io3_di 0.01fF
C7223 raven_soc_0|gpio_outenb<4> raven_soc_0|ext_clk 0.01fF
C7224 BU_3VX2_31|A vdd 0.86fF
C7225 BU_3VX2_26|A raven_soc_0|flash_io2_do 0.01fF
C7226 raven_soc_0|gpio_pullup<0> BU_3VX2_27|Q 0.03fF
C7227 VDD raven_padframe_0|APR00DF_2|GNDO 0.07fF
C7228 raven_soc_0|gpio_pulldown<2> BU_3VX2_28|Q 0.01fF
C7229 raven_soc_0|gpio_out<10> raven_soc_0|gpio_outenb<8> 5.31fF
C7230 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<6> 0.08fF
C7231 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<10> 21.96fF
C7232 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<31> 181.10fF
C7233 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<7> 2.63fF
C7234 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<24> 0.01fF
C7235 BU_3VX2_32|Q BU_3VX2_11|Q 8.91fF
C7236 BU_3VX2_37|Q BU_3VX2_36|Q 0.75fF
C7237 BU_3VX2_70|Q BU_3VX2_4|Q 1.46fF
C7238 raven_padframe_0|ICF_2|GNDR raven_padframe_0|ICF_2|GNDO 0.81fF
C7239 raven_padframe_0|BBC4F_2|GNDR raven_padframe_0|BBC4F_2|VDDO 0.09fF
C7240 raven_padframe_0|BT4F_0|GNDR raven_padframe_0|BT4F_0|GNDO 0.81fF
C7241 raven_padframe_0|BBCUD4F_8|GNDR raven_padframe_0|BBCUD4F_8|VDDO 0.09fF
C7242 BU_3VX2_24|A raven_soc_0|flash_io0_di 0.01fF
C7243 raven_soc_0|gpio_out<0> raven_soc_0|flash_io3_do 5.50fF
C7244 raven_soc_0|gpio_outenb<1> LS_3VX2_3|A 0.81fF
C7245 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<12> 0.01fF
C7246 raven_padframe_0|BBC4F_0|VDDR raven_padframe_0|BBC4F_0|GNDO 0.13fF
C7247 BU_3VX2_67|A BU_3VX2_66|Q 0.16fF
C7248 LS_3VX2_11|Q LS_3VX2_22|A 0.01fF
C7249 raven_soc_0|gpio_pullup<2> BU_3VX2_23|Q 0.01fF
C7250 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<10> 0.94fF
C7251 VDD raven_padframe_0|VDDORPADF_0|GNDO 0.07fF
C7252 BU_3VX2_11|A raven_soc_0|flash_io2_do 0.01fF
C7253 VDD raven_padframe_0|BBCUD4F_11|GNDR 0.16fF
C7254 raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<15> 13.44fF
C7255 BU_3VX2_36|A BU_3VX2_32|Q 0.02fF
C7256 BU_3VX2_0|Q raven_soc_0|ram_rdata<23> 0.02fF
C7257 BU_3VX2_10|A BU_3VX2_21|A 1.16fF
C7258 VDD raven_padframe_0|BBC4F_3|VDDR 0.71fF
C7259 BU_3VX2_63|A BU_3VX2_17|A 0.01fF
C7260 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_out<4> 1.20fF
C7261 BU_3VX2_18|A BU_3VX2_13|A 3.87fF
C7262 BU_3VX2_40|A BU_3VX2_31|A 0.02fF
C7263 BU_3VX2_1|A BU_3VX2_33|A 0.28fF
C7264 BU_3VX2_31|A raven_soc_0|gpio_in<2> 0.01fF
C7265 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<14> 2.25fF
C7266 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<8> 0.02fF
C7267 raven_soc_0|gpio_out<9> raven_soc_0|gpio_outenb<8> 11.38fF
C7268 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<14> 12.13fF
C7269 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<5> 0.01fF
C7270 raven_soc_0|gpio_out<7> BU_3VX2_71|Q 0.01fF
C7271 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<8> 0.01fF
C7272 raven_soc_0|gpio_out<11> raven_soc_0|gpio_outenb<13> 7.57fF
C7273 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<1> 9.23fF
C7274 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<9> 0.01fF
C7275 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<8> 0.01fF
C7276 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<5> 4.48fF
C7277 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<13> 0.44fF
C7278 BU_3VX2_13|Q BU_3VX2_8|Q 10.99fF
C7279 BU_3VX2_38|Q BU_3VX2_17|Q 46.53fF
C7280 raven_soc_0|ram_wdata<1> raven_soc_0|ram_rdata<13> 0.76fF
C7281 BU_3VX2_13|Q BU_3VX2_21|Q 10.69fF
C7282 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<19> 9.92fF
C7283 BU_3VX2_66|Q BU_3VX2_10|Q 0.02fF
C7284 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<25> 20.81fF
C7285 BU_3VX2_2|Q BU_3VX2_66|Q 1.86fF
C7286 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<22> 15.84fF
C7287 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<26> 0.03fF
C7288 BU_3VX2_1|Q BU_3VX2_64|Q 0.77fF
C7289 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<29> 7.04fF
C7290 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<1> 0.01fF
C7291 LS_3VX2_18|A AMUX4_3V_4|SEL[1] 1.02fF
C7292 BU_3VX2_10|Q BU_3VX2_20|Q 7.66fF
C7293 BU_3VX2_67|Q BU_3VX2_17|Q 0.11fF
C7294 VDD3V3 BU_3VX2_29|Q 1.86fF
C7295 raven_soc_0|ext_clk apllc03_1v8_0|CLK 97.89fF
C7296 LS_3VX2_16|Q vdd 0.40fF
C7297 raven_soc_0|gpio_in<14> BU_3VX2_24|Q 0.01fF
C7298 raven_soc_0|gpio_in<12> BU_3VX2_26|Q 0.01fF
C7299 LS_3VX2_20|Q BU_3VX2_45|Q 0.30fF
C7300 raven_soc_0|gpio_in<9> BU_3VX2_25|Q 0.01fF
C7301 BU_3VX2_21|A BU_3VX2_0|A 0.20fF
C7302 raven_padframe_0|BBC4F_3|VDDR LOGIC0_3V_4|Q 0.01fF
C7303 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_in<4> 1.02fF
C7304 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<10> 0.31fF
C7305 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<4> 0.41fF
C7306 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<4> 0.01fF
C7307 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<11> 0.01fF
C7308 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<15> 0.02fF
C7309 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<0> 0.01fF
C7310 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<13> 0.07fF
C7311 raven_soc_0|gpio_out<8> vdd 0.21fF
C7312 BU_3VX2_3|Q vdd 1.55fF
C7313 raven_soc_0|ram_rdata<17> apllc03_1v8_0|CLK 0.01fF
C7314 LS_3VX2_13|Q vdd 0.16fF
C7315 BU_3VX2_31|A raven_soc_0|gpio_in<11> 0.01fF
C7316 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<6> 1.14fF
C7317 LS_3VX2_3|A raven_soc_0|gpio_pulldown<3> 0.37fF
C7318 BU_3VX2_0|Q raven_soc_0|ram_wdata<21> 0.02fF
C7319 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<16> 6.86fF
C7320 BU_3VX2_41|A BU_3VX2_46|Q 0.15fF
C7321 raven_padframe_0|FILLER20F_0|GNDR raven_padframe_0|FILLER20F_0|VDDO 0.09fF
C7322 raven_padframe_0|APR00DF_6|VDDR raven_padframe_0|APR00DF_6|GNDR 0.68fF
C7323 acmpc01_3v3_0|IBN acsoc01_3v3_0|CS2_200N 0.04fF
C7324 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<5> 0.49fF
C7325 BU_3VX2_32|A BU_3VX2_68|A 0.54fF
C7326 BU_3VX2_7|A BU_3VX2_38|A 1.05fF
C7327 LS_3VX2_18|Q vdd 0.33fF
C7328 BU_3VX2_63|A BU_3VX2_12|A 0.01fF
C7329 BU_3VX2_23|A raven_soc_0|flash_io2_oeb 2.84fF
C7330 BU_3VX2_22|A vdd 0.06fF
C7331 BU_3VX2_16|A raven_soc_0|flash_io0_di 0.11fF
C7332 raven_padframe_0|ICFC_2|VDDR raven_padframe_0|ICFC_2|VDDO 0.06fF
C7333 raven_padframe_0|POWERCUTVDD3FC_1|VDDR raven_padframe_0|POWERCUTVDD3FC_1|GNDR 0.64fF
C7334 LS_3VX2_11|A LS_3VX2_27|A 6.01fF
C7335 LS_3VX2_8|A LS_3VX2_19|A 0.01fF
C7336 BU_3VX2_31|A raven_soc_0|gpio_outenb<9> 0.01fF
C7337 LS_3VX2_8|A BU_3VX2_52|Q 8.19fF
C7338 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<8> 0.01fF
C7339 BU_3VX2_29|A raven_soc_0|flash_io0_di 0.01fF
C7340 IN_3VX2_1|A BU_3VX2_27|Q 44.80fF
C7341 raven_padframe_0|BBCUD4F_8|VDDR raven_padframe_0|BBCUD4F_8|GNDR 0.68fF
C7342 raven_soc_0|gpio_out<6> vdd 0.19fF
C7343 raven_soc_0|gpio_outenb<11> BU_3VX2_28|Q 0.01fF
C7344 raven_soc_0|gpio_outenb<10> apllc03_1v8_0|CLK 0.01fF
C7345 raven_soc_0|gpio_outenb<15> BU_3VX2_24|Q 0.01fF
C7346 raven_soc_0|gpio_outenb<14> BU_3VX2_23|Q 0.01fF
C7347 raven_padframe_0|BBCUD4F_4|VDDR raven_padframe_0|BBCUD4F_4|GNDR 0.68fF
C7348 raven_soc_0|gpio_in<1> LS_3VX2_3|A 0.39fF
C7349 BU_3VX2_23|A BU_3VX2_6|A 0.01fF
C7350 BU_3VX2_19|A BU_3VX2_4|A 0.01fF
C7351 BU_3VX2_65|A BU_3VX2_70|A 2.50fF
C7352 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<14> 1.27fF
C7353 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<9> 0.01fF
C7354 BU_3VX2_37|A raven_soc_0|flash_io0_di 0.01fF
C7355 LS_3VX2_3|A raven_soc_0|gpio_outenb<5> 0.01fF
C7356 BU_3VX2_35|A raven_soc_0|flash_clk 0.01fF
C7357 BU_3VX2_0|Q raven_soc_0|gpio_pullup<4> 0.01fF
C7358 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<11> 12.73fF
C7359 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<11> 14.54fF
C7360 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<8> 0.02fF
C7361 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<14> 0.01fF
C7362 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<23> 0.01fF
C7363 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<10> 7.09fF
C7364 raven_soc_0|gpio_in<6> raven_soc_0|gpio_in<15> 6.23fF
C7365 AMUX4_3V_3|SEL[1] BU_3VX2_68|Q 0.26fF
C7366 raven_soc_0|gpio_in<14> raven_soc_0|gpio_out<15> 50.89fF
C7367 BU_3VX2_24|A BU_3VX2_5|A 0.01fF
C7368 LS_3VX2_16|Q BU_3VX2_62|A 1.87fF
C7369 raven_soc_0|flash_io2_do VDD3V3 12.34fF
C7370 LOGIC0_3V_1|Q BU_3VX2_33|A 3.61fF
C7371 BU_3VX2_9|A BU_3VX2_35|A 0.62fF
C7372 LS_3VX2_11|A LS_3VX2_10|Q 0.16fF
C7373 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<1> 8.25fF
C7374 raven_padframe_0|FILLER20FC_0|VDD3 BU_3VX2_33|A 0.01fF
C7375 BU_3VX2_71|A BU_3VX2_13|A 0.01fF
C7376 BU_3VX2_20|A raven_soc_0|flash_csb 1.74fF
C7377 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<4> 1.03fF
C7378 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<9> 0.01fF
C7379 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<9> 1.29fF
C7380 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<6> 0.02fF
C7381 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<12> 0.33fF
C7382 markings_0|efabless_logo_0|m1_3600_n10650# markings_0|efabless_logo_0|m1_4500_n11550# 0.37fF
C7383 markings_0|efabless_logo_0|m1_2700_n10050# markings_0|efabless_logo_0|m2_3000_n6450# 0.01fF
C7384 LS_3VX2_7|A LS_3VX2_20|A 5.29fF
C7385 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<11> 1.37fF
C7386 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<25> 16.55fF
C7387 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<2> 0.01fF
C7388 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<14> 0.30fF
C7389 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<12> 27.12fF
C7390 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<15> 0.54fF
C7391 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<14> 0.01fF
C7392 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<19> 0.12fF
C7393 BU_3VX2_71|Q BU_3VX2_40|Q 37.23fF
C7394 raven_soc_0|gpio_out<14> raven_soc_0|gpio_pullup<5> 0.02fF
C7395 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<15> 0.01fF
C7396 raven_soc_0|gpio_outenb<8> raven_soc_0|ext_clk 0.01fF
C7397 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_out<15> 0.02fF
C7398 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<7> 0.01fF
C7399 raven_soc_0|ram_rdata<18> vdd 0.36fF
C7400 BU_3VX2_62|Q BU_3VX2_53|Q 12.86fF
C7401 LS_3VX2_12|A LS_3VX2_13|A 55.77fF
C7402 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<11> 0.01fF
C7403 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<8> 0.94fF
C7404 LS_3VX2_9|A BU_3VX2_57|Q 11.17fF
C7405 VDD raven_padframe_0|CORNERESDF_3|GNDO 0.07fF
C7406 LS_3VX2_5|A BU_3VX2_53|Q 17.86fF
C7407 BU_3VX2_0|Q BU_3VX2_2|Q 0.01fF
C7408 LS_3VX2_4|A LS_3VX2_19|A 0.49fF
C7409 analog_out AMUX4_3V_4|AIN2 11.91fF
C7410 raven_soc_0|gpio_pullup<0> BU_3VX2_25|Q 0.01fF
C7411 LS_3VX2_4|A BU_3VX2_52|Q 34.20fF
C7412 raven_soc_0|gpio_pulldown<2> vdd 0.20fF
C7413 BU_3VX2_0|Q BU_3VX2_10|Q 0.01fF
C7414 VDD raven_padframe_0|CORNERESDF_1|GNDO 0.07fF
C7415 raven_soc_0|gpio_out<8> raven_soc_0|gpio_outenb<9> 9.87fF
C7416 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<5> 0.08fF
C7417 BU_3VX2_3|Q BU_3VX2_70|Q 4.23fF
C7418 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<6> 2.17fF
C7419 raven_soc_0|ram_rdata<24> raven_soc_0|ram_addr<2> 5.34fF
C7420 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<10> 3.05fF
C7421 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<9> 7.96fF
C7422 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<31> 1.35fF
C7423 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<20> 0.06fF
C7424 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<6> 0.01fF
C7425 raven_soc_0|ram_wdata<23> raven_soc_0|ram_addr<4> 0.01fF
C7426 LS_3VX2_27|A LS_3VX2_21|A 164.68fF
C7427 raven_padframe_0|axtoc02_3v3_0|GNDR raven_padframe_0|axtoc02_3v3_0|VDDO 0.14fF
C7428 LS_3VX2_3|Q raven_soc_0|flash_io0_di 0.01fF
C7429 BU_3VX2_21|A vdd 0.06fF
C7430 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<13> 10.97fF
C7431 raven_padframe_0|GNDORPADF_5|VDDR raven_padframe_0|GNDORPADF_5|GNDOR 0.81fF
C7432 IN_3VX2_1|A raven_soc_0|flash_io2_oeb 19.97fF
C7433 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<15> 0.39fF
C7434 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<15> 312.91fF
C7435 LOGIC0_3V_4|Q raven_padframe_0|BBC4F_1|PO 0.04fF
C7436 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<8> 3.59fF
C7437 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<11> 0.16fF
C7438 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<15> 0.02fF
C7439 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<6> 0.13fF
C7440 BU_3VX2_0|Q raven_soc_0|flash_clk 0.21fF
C7441 BU_3VX2_33|A BU_3VX2_1|Q 0.03fF
C7442 BU_3VX2_6|A IN_3VX2_1|A 0.01fF
C7443 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<2> 91.87fF
C7444 AMUX4_3V_0|AIN1 BU_3VX2_51|A 0.02fF
C7445 LOGIC0_3V_4|Q raven_soc_0|flash_io0_di 0.10fF
C7446 LS_3VX2_8|A BU_3VX2_58|Q 0.01fF
C7447 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<8> 6.44fF
C7448 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<14> 10.95fF
C7449 raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<10> 1.46fF
C7450 raven_soc_0|gpio_outenb<7> BU_3VX2_71|Q 0.01fF
C7451 raven_soc_0|gpio_out<6> raven_soc_0|gpio_outenb<9> 0.01fF
C7452 raven_soc_0|gpio_out<1> VDD3V3 1.61fF
C7453 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<5> 0.01fF
C7454 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pullup<13> 0.01fF
C7455 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pullup<14> 0.01fF
C7456 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<27> 0.08fF
C7457 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<29> 0.16fF
C7458 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<26> 0.35fF
C7459 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<25> 0.13fF
C7460 BU_3VX2_19|Q BU_3VX2_13|Q 5.98fF
C7461 BU_3VX2_13|Q BU_3VX2_18|Q 11.80fF
C7462 BU_3VX2_21|Q BU_3VX2_69|Q 2.52fF
C7463 BU_3VX2_2|Q BU_3VX2_30|Q 0.24fF
C7464 BU_3VX2_16|Q BU_3VX2_10|Q 6.28fF
C7465 BU_3VX2_12|Q BU_3VX2_9|Q 14.46fF
C7466 BU_3VX2_6|Q BU_3VX2_22|Q 4.11fF
C7467 BU_3VX2_15|Q BU_3VX2_12|Q 13.57fF
C7468 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<17> 0.23fF
C7469 BU_3VX2_16|Q BU_3VX2_2|Q 0.49fF
C7470 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<19> 7.26fF
C7471 raven_soc_0|ram_wdata<15> raven_soc_0|ram_rdata<2> 0.01fF
C7472 BU_3VX2_66|Q BU_3VX2_33|Q 0.53fF
C7473 BU_3VX2_30|Q BU_3VX2_10|Q 2.84fF
C7474 BU_3VX2_7|Q BU_3VX2_22|Q 5.65fF
C7475 BU_3VX2_69|Q BU_3VX2_8|Q 0.44fF
C7476 AMUX4_3V_0|SEL[1] BU_3VX2_42|Q 7.33fF
C7477 BU_3VX2_53|A vdd 0.07fF
C7478 BU_3VX2_43|A BU_3VX2_44|Q 0.03fF
C7479 BU_3VX2_42|Q BU_3VX2_51|Q 58.12fF
C7480 LOGIC1_3V_1|Q LOGIC1_3V_0|Q 0.58fF
C7481 raven_padframe_0|POWERCUTVDD3FC_1|VDDO raven_padframe_0|POWERCUTVDD3FC_1|GNDO 2.22fF
C7482 BU_3VX2_5|A BU_3VX2_16|A 0.96fF
C7483 raven_soc_0|gpio_pullup<2> BU_3VX2_31|A 0.04fF
C7484 BU_3VX2_23|A BU_3VX2_27|A 10.04fF
C7485 LS_3VX2_12|A raven_soc_0|ser_rx 0.01fF
C7486 BU_3VX2_5|A BU_3VX2_29|A 0.01fF
C7487 BU_3VX2_35|A BU_3VX2_28|A 0.01fF
C7488 raven_padframe_0|aregc01_3v3_1|m4_0_31172# raven_padframe_0|aregc01_3v3_1|m4_0_30653# 0.09fF
C7489 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<10> 0.01fF
C7490 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<10> 7.97fF
C7491 BU_3VX2_1|Q raven_soc_0|flash_io3_do 0.01fF
C7492 raven_soc_0|gpio_pulldown<6> vdd 0.36fF
C7493 AMUX4_3V_3|SEL[1] BU_3VX2_24|Q 1.49fF
C7494 raven_soc_0|irq_pin BU_3VX2_59|Q 0.01fF
C7495 raven_soc_0|ram_wdata<22> apllc03_1v8_0|CLK 0.01fF
C7496 BU_3VX2_37|A BU_3VX2_5|A 2.21fF
C7497 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<12> 0.03fF
C7498 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<13> 0.01fF
C7499 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<13> 1.61fF
C7500 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<11> 0.34fF
C7501 raven_soc_0|gpio_outenb<3> BU_3VX2_40|Q 0.77fF
C7502 raven_padframe_0|APR00DF_0|VDDR raven_padframe_0|APR00DF_0|GNDO 0.13fF
C7503 raven_soc_0|flash_io0_di raven_soc_0|flash_io1_oeb 16.59fF
C7504 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<1> 0.01fF
C7505 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<16> 0.18fF
C7506 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<15> 0.05fF
C7507 raven_soc_0|ram_rdata<9> raven_soc_0|ram_addr<0> 0.03fF
C7508 raven_soc_0|flash_io3_di raven_soc_0|flash_clk 15.10fF
C7509 BU_3VX2_47|A BU_3VX2_45|Q 0.02fF
C7510 raven_padframe_0|ICFC_0|VDDO raven_padframe_0|ICFC_0|GNDO 2.28fF
C7511 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<6> 0.30fF
C7512 BU_3VX2_24|A BU_3VX2_24|Q 0.08fF
C7513 BU_3VX2_9|A raven_soc_0|flash_io3_di 0.01fF
C7514 LS_3VX2_9|A LS_3VX2_16|A 0.08fF
C7515 BU_3VX2_7|A BU_3VX2_4|Q 0.02fF
C7516 BU_3VX2_19|A raven_soc_0|flash_io0_oeb 0.01fF
C7517 LS_3VX2_8|A LS_3VX2_22|A 23.30fF
C7518 raven_padframe_0|BT4FC_0|VDDR raven_padframe_0|BT4FC_0|GNDR 0.68fF
C7519 LS_3VX2_7|A BU_3VX2_47|Q 0.26fF
C7520 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<9> 0.60fF
C7521 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<6> 0.01fF
C7522 IN_3VX2_1|A BU_3VX2_25|Q 31.64fF
C7523 LS_3VX2_4|A BU_3VX2_58|Q 9.85fF
C7524 raven_soc_0|gpio_pullup<10> apllc03_1v8_0|CLK 0.01fF
C7525 raven_soc_0|gpio_outenb<11> vdd 0.22fF
C7526 raven_soc_0|gpio_pullup<8> BU_3VX2_29|Q 0.01fF
C7527 raven_soc_0|gpio_pullup<11> BU_3VX2_28|Q 0.01fF
C7528 raven_soc_0|gpio_pullup<15> BU_3VX2_23|Q 0.01fF
C7529 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<15> 0.01fF
C7530 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<9> 0.94fF
C7531 LS_3VX2_3|A raven_soc_0|gpio_pullup<7> 0.01fF
C7532 BU_3VX2_25|A raven_soc_0|flash_io2_oeb 2.97fF
C7533 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<11> 26.64fF
C7534 LS_3VX2_6|A BU_3VX2_59|Q 5.78fF
C7535 BU_3VX2_63|Q raven_soc_0|flash_io1_oeb 0.22fF
C7536 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<6> 1.07fF
C7537 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<7> 4.92fF
C7538 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<8> 15.92fF
C7539 raven_soc_0|ext_clk raven_soc_0|gpio_in<15> 0.01fF
C7540 BU_3VX2_54|A LS_3VX2_17|Q 0.11fF
C7541 BU_3VX2_56|A LS_3VX2_15|Q 0.22fF
C7542 BU_3VX2_58|A BU_3VX2_60|A 2.18fF
C7543 BU_3VX2_55|A LS_3VX2_16|Q 0.15fF
C7544 BU_3VX2_57|A BU_3VX2_61|A 0.60fF
C7545 BU_3VX2_53|A BU_3VX2_62|A 0.13fF
C7546 BU_3VX2_24|A BU_3VX2_13|A 1.91fF
C7547 BU_3VX2_43|A vdd 0.06fF
C7548 BU_3VX2_6|A BU_3VX2_25|A 0.01fF
C7549 BU_3VX2_5|A LS_3VX2_3|Q 0.64fF
C7550 IN_3VX2_1|A BU_3VX2_27|A 19.21fF
C7551 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<1> 20.84fF
C7552 raven_padframe_0|aregc01_3v3_0|m4_0_31172# raven_padframe_0|aregc01_3v3_0|m4_0_30133# 0.02fF
C7553 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<7> 1.82fF
C7554 BU_3VX2_31|A raven_soc_0|gpio_outenb<14> 0.01fF
C7555 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<11> 0.01fF
C7556 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<0> 7.02fF
C7557 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<9> 0.01fF
C7558 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<20> 1.31fF
C7559 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<14> 0.30fF
C7560 raven_soc_0|gpio_pullup<14> BU_3VX2_40|Q 0.02fF
C7561 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<6> 9.02fF
C7562 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<11> 0.02fF
C7563 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<12> 14.67fF
C7564 raven_soc_0|flash_clk raven_soc_0|irq_pin 0.06fF
C7565 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<0> 0.05fF
C7566 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<1> 0.01fF
C7567 BU_3VX2_13|Q BU_3VX2_27|Q 2.15fF
C7568 LS_3VX2_19|A vdd 3.24fF
C7569 BU_3VX2_21|Q BU_3VX2_29|Q 6.12fF
C7570 BU_3VX2_52|Q vdd 1.77fF
C7571 LS_3VX2_20|Q LS_3VX2_21|A 0.19fF
C7572 BU_3VX2_8|Q BU_3VX2_29|Q 0.01fF
C7573 LOGIC0_3V_4|Q raven_soc_0|gpio_out<2> 0.74fF
C7574 IN_3VX2_1|Q LS_3VX2_20|A 0.01fF
C7575 raven_padframe_0|FILLER20FC_0|VDDR raven_padframe_0|FILLER20FC_0|GNDO 0.13fF
C7576 LS_3VX2_4|A LS_3VX2_22|A 7.94fF
C7577 AMUX4_3V_4|AIN1 AMUX4_3V_4|AIN2 57.83fF
C7578 BU_3VX2_0|Q BU_3VX2_33|Q 0.01fF
C7579 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_out<10> 0.02fF
C7580 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_outenb<13> 0.02fF
C7581 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_outenb<9> 1.94fF
C7582 AMUX4_3V_3|SEL[1] LS_3VX2_23|A 8.95fF
C7583 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<8> 0.37fF
C7584 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<4> 0.85fF
C7585 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<30> 0.51fF
C7586 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<24> 14.37fF
C7587 raven_soc_0|ram_rdata<22> raven_soc_0|ram_addr<3> 4.01fF
C7588 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<23> 0.01fF
C7589 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<10> 12.66fF
C7590 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<5> 0.01fF
C7591 BU_3VX2_63|A raven_soc_0|flash_clk 0.01fF
C7592 VDD raven_padframe_0|BBCUD4F_15|GNDO 0.07fF
C7593 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<14> 0.03fF
C7594 BU_3VX2_12|A BU_3VX2_11|Q 0.16fF
C7595 BU_3VX2_28|A raven_soc_0|flash_io3_di 0.01fF
C7596 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<11> 141.28fF
C7597 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<9> 2.12fF
C7598 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<14> 0.17fF
C7599 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<6> 0.07fF
C7600 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<12> 0.03fF
C7601 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<15> 0.17fF
C7602 adc_low vdd 1.61fF
C7603 raven_soc_0|gpio_out<13> raven_soc_0|ext_clk 0.01fF
C7604 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pullup<5> 0.02fF
C7605 raven_soc_0|gpio_out<11> VDD3V3 0.07fF
C7606 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<23> 2.74fF
C7607 BU_3VX2_9|A BU_3VX2_63|A 0.02fF
C7608 BU_3VX2_7|A BU_3VX2_31|A 0.01fF
C7609 BU_3VX2_68|A BU_3VX2_64|A 3.31fF
C7610 BU_3VX2_5|A raven_soc_0|flash_io1_oeb 0.01fF
C7611 BU_3VX2_25|A BU_3VX2_25|Q 0.08fF
C7612 LS_3VX2_8|A BU_3VX2_60|Q 0.02fF
C7613 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<3> 0.01fF
C7614 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<6> 0.01fF
C7615 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<8> 3.60fF
C7616 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pullup<14> 0.02fF
C7617 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<10> 1.41fF
C7618 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<8> 0.10fF
C7619 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<9> 7.36fF
C7620 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<14> 18.25fF
C7621 raven_soc_0|gpio_pullup<9> BU_3VX2_71|Q 0.01fF
C7622 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pullup<6> 2.05fF
C7623 raven_soc_0|gpio_pulldown<8> BU_3VX2_28|Q 0.01fF
C7624 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<15> 103.43fF
C7625 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<12> 1.15fF
C7626 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<25> 0.15fF
C7627 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<2> 0.01fF
C7628 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<17> 2.48fF
C7629 BU_3VX2_15|Q BU_3VX2_5|Q 5.46fF
C7630 BU_3VX2_38|Q BU_3VX2_68|Q 0.86fF
C7631 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<13> 0.50fF
C7632 raven_soc_0|ram_wdata<8> raven_soc_0|ram_rdata<25> 0.56fF
C7633 raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<15> 2.08fF
C7634 BU_3VX2_12|Q BU_3VX2_64|Q 0.39fF
C7635 BU_3VX2_19|Q BU_3VX2_69|Q 3.05fF
C7636 BU_3VX2_68|Q BU_3VX2_67|Q 40.09fF
C7637 BU_3VX2_69|Q BU_3VX2_18|Q 1.38fF
C7638 VDD3V3 AMUX4_3V_4|AIN2 19.66fF
C7639 BU_3VX2_31|Q BU_3VX2_7|Q 0.33fF
C7640 BU_3VX2_5|Q BU_3VX2_9|Q 10.07fF
C7641 BU_3VX2_73|Q BU_3VX2_55|Q 0.01fF
C7642 BU_3VX2_42|Q BU_3VX2_49|Q 28.11fF
C7643 BU_3VX2_44|A BU_3VX2_43|Q 0.14fF
C7644 raven_padframe_0|CORNERESDF_3|VDDR raven_padframe_0|CORNERESDF_3|VDDO 0.06fF
C7645 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<2> 92.25fF
C7646 BU_3VX2_16|A BU_3VX2_13|A 7.16fF
C7647 BU_3VX2_35|A LS_3VX2_3|A 0.55fF
C7648 BU_3VX2_13|A BU_3VX2_29|A 0.01fF
C7649 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<3> 4.81fF
C7650 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<4> 1.95fF
C7651 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<12> 0.93fF
C7652 raven_soc_0|gpio_pulldown<15> LS_3VX2_3|A 0.01fF
C7653 raven_soc_0|gpio_pulldown<13> BU_3VX2_63|Q 0.01fF
C7654 raven_padframe_0|CORNERESDF_1|GNDR raven_padframe_0|CORNERESDF_1|VDDO 0.09fF
C7655 raven_soc_0|flash_io3_di BU_3VX2_33|Q 0.01fF
C7656 raven_soc_0|irq_pin BU_3VX2_61|Q 0.01fF
C7657 raven_soc_0|ram_rdata<27> apllc03_1v8_0|CLK 0.01fF
C7658 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<0> 29.09fF
C7659 BU_3VX2_37|A BU_3VX2_13|A 1.16fF
C7660 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<12> 0.25fF
C7661 BU_3VX2_25|A BU_3VX2_27|A 20.59fF
C7662 LS_3VX2_6|A AMUX2_3V_0|SEL 12.81fF
C7663 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<5> 0.01fF
C7664 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<12> 168.23fF
C7665 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<13> 0.65fF
C7666 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<9> 1.15fF
C7667 raven_soc_0|gpio_pullup<1> BU_3VX2_63|Q 0.04fF
C7668 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<6> 0.01fF
C7669 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<15> 0.01fF
C7670 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<11> 0.02fF
C7671 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<14> 0.01fF
C7672 BU_3VX2_18|A raven_soc_0|ext_clk 0.01fF
C7673 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<31> 7.03fF
C7674 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<1> 0.05fF
C7675 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<13> 0.03fF
C7676 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<25> 168.38fF
C7677 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io2_di 37.96fF
C7678 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<15> 10.95fF
C7679 raven_soc_0|ram_rdata<14> raven_soc_0|ram_addr<0> 0.41fF
C7680 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<16> 0.06fF
C7681 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<17> 1.87fF
C7682 BU_3VX2_36|Q BU_3VX2_17|Q 1.56fF
C7683 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<21> 0.07fF
C7684 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<31> 0.01fF
C7685 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<27> 0.01fF
C7686 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<29> 3.05fF
C7687 BU_3VX2_58|Q vdd 2.07fF
C7688 raven_padframe_0|FILLER20F_2|VDDR raven_padframe_0|FILLER20F_2|VDDO 0.06fF
C7689 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<8> 0.01fF
C7690 BU_3VX2_2|A raven_soc_0|flash_io2_di 0.02fF
C7691 BU_3VX2_19|A raven_soc_0|flash_io2_do 0.01fF
C7692 LS_3VX2_11|A BU_3VX2_53|Q 13.17fF
C7693 BU_3VX2_4|A raven_soc_0|flash_io2_oeb 0.01fF
C7694 raven_padframe_0|FILLER20FC_0|VDD3 raven_padframe_0|FILLER20FC_0|GNDR 0.16fF
C7695 raven_padframe_0|GNDORPADF_3|VDDR raven_padframe_0|GNDORPADF_3|VDDO 0.06fF
C7696 IN_3VX2_1|A AMUX4_3V_0|SEL[1] 17.94fF
C7697 LS_3VX2_4|A BU_3VX2_60|Q 7.84fF
C7698 IN_3VX2_1|A BU_3VX2_51|Q 0.01fF
C7699 raven_soc_0|gpio_pullup<11> vdd 0.39fF
C7700 AMUX2_3V_0|AOUT vdd 0.03fF
C7701 raven_soc_0|gpio_pulldown<4> apllc03_1v8_0|CLK 0.01fF
C7702 BU_3VX2_6|A BU_3VX2_4|A 7.60fF
C7703 BU_3VX2_68|A BU_3VX2_66|A 8.45fF
C7704 BU_3VX2_63|A BU_3VX2_28|A 0.01fF
C7705 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<6> 0.01fF
C7706 XSPRAM_1024X32_M8P_0|RDY BU_3VX2_0|Q 0.06fF
C7707 LS_3VX2_12|A AMUX4_3V_1|SEL[0] 9.70fF
C7708 LS_3VX2_3|A BU_3VX2_0|Q 55.88fF
C7709 BU_3VX2_35|A raven_soc_0|flash_io1_do 0.07fF
C7710 AMUX4_3V_4|AOUT raven_soc_0|flash_io2_oeb 0.47fF
C7711 IN_3VX2_1|Q BU_3VX2_47|Q 0.68fF
C7712 BU_3VX2_14|A raven_soc_0|flash_io3_di 0.01fF
C7713 VDD raven_padframe_0|BBCUD4F_6|GNDO 0.07fF
C7714 LS_3VX2_6|A BU_3VX2_61|Q 0.01fF
C7715 raven_soc_0|ext_clk raven_soc_0|gpio_in<14> 0.01fF
C7716 BU_3VX2_40|Q raven_soc_0|gpio_in<9> 0.01fF
C7717 raven_soc_0|gpio_in<12> VDD3V3 0.07fF
C7718 BU_3VX2_52|A BU_3VX2_56|A 1.39fF
C7719 BU_3VX2_53|A BU_3VX2_55|A 4.05fF
C7720 VDD3V3 BU_3VX2_58|A 0.05fF
C7721 BU_3VX2_22|A BU_3VX2_7|A 0.67fF
C7722 AMUX4_3V_3|AOUT AMUX4_3V_4|AIN1 0.02fF
C7723 LS_3VX2_3|Q BU_3VX2_13|A 0.01fF
C7724 BU_3VX2_17|A BU_3VX2_26|A 2.38fF
C7725 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<9> 3.30fF
C7726 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<12> 0.01fF
C7727 raven_soc_0|gpio_pulldown<0> LS_3VX2_3|A 0.01fF
C7728 BU_3VX2_31|A raven_soc_0|gpio_pullup<15> 0.01fF
C7729 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<11> 0.01fF
C7730 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<2> 0.01fF
C7731 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<10> 0.01fF
C7732 markings_0|efabless_logo_0|m1_7500_n3450# markings_0|efabless_logo_0|m1_8400_n4650# 0.19fF
C7733 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<20> 0.46fF
C7734 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<0> 0.01fF
C7735 raven_soc_0|gpio_pullup<6> raven_soc_0|ext_clk 0.04fF
C7736 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<8> 8.93fF
C7737 LS_3VX2_22|A vdd 4.33fF
C7738 BU_3VX2_13|Q BU_3VX2_25|Q 3.37fF
C7739 BU_3VX2_38|Q BU_3VX2_24|Q 9.37fF
C7740 BU_3VX2_2|Q BU_3VX2_26|Q 0.03fF
C7741 BU_3VX2_6|Q apllc03_1v8_0|CLK 0.01fF
C7742 BU_3VX2_15|Q BU_3VX2_28|Q 2.70fF
C7743 BU_3VX2_19|Q BU_3VX2_29|Q 3.40fF
C7744 BU_3VX2_67|Q BU_3VX2_24|Q 0.84fF
C7745 BU_3VX2_22|Q BU_3VX2_23|Q 66.04fF
C7746 BU_3VX2_18|Q BU_3VX2_29|Q 3.92fF
C7747 BU_3VX2_69|Q BU_3VX2_27|Q 0.34fF
C7748 BU_3VX2_9|Q BU_3VX2_28|Q 0.43fF
C7749 BU_3VX2_10|Q BU_3VX2_26|Q 0.02fF
C7750 BU_3VX2_7|Q apllc03_1v8_0|CLK 0.01fF
C7751 LS_3VX2_20|Q LS_3VX2_27|A 0.01fF
C7752 raven_padframe_0|BT4FC_0|VDD3 LOGIC0_3V_4|Q 0.04fF
C7753 BU_3VX2_17|A BU_3VX2_11|A 3.05fF
C7754 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<11> 0.01fF
C7755 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<1> 106.82fF
C7756 BU_3VX2_33|A LOGIC0_3V_2|Q 1.33fF
C7757 BU_3VX2_10|A BU_3VX2_9|Q 0.16fF
C7758 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<10> 0.01fF
C7759 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pullup<13> 0.02fF
C7760 raven_soc_0|ram_rdata<17> raven_soc_0|ram_rdata<15> 33.69fF
C7761 raven_soc_0|flash_io2_di apllc03_1v8_0|CLK 23.77fF
C7762 raven_soc_0|ram_rdata<20> vdd 0.61fF
C7763 raven_soc_0|flash_io1_oeb BU_3VX2_24|Q 0.01fF
C7764 raven_soc_0|flash_io0_oeb BU_3VX2_27|Q 0.01fF
C7765 raven_soc_0|flash_clk BU_3VX2_26|Q 0.01fF
C7766 BU_3VX2_46|Q BU_3VX2_72|Q 1.44fF
C7767 raven_padframe_0|FILLER01F_1|VDDO raven_padframe_0|FILLER01F_1|GNDO 2.28fF
C7768 raven_padframe_0|FILLER50F_0|GNDR raven_padframe_0|FILLER50F_0|VDDO 0.09fF
C7769 raven_padframe_0|aregc01_3v3_1|GNDR raven_padframe_0|aregc01_3v3_1|VDDO 0.07fF
C7770 markings_0|date_0|_alphabet_2_0|m2_0_0# markings_0|manufacturer_0|_alphabet_L_0|m2_0_0# 0.11fF
C7771 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<13> 0.78fF
C7772 VDD raven_soc_0|gpio_out<15> 0.01fF
C7773 AMUX4_3V_3|AOUT VDD3V3 5.77fF
C7774 BU_3VX2_1|A BU_3VX2_1|Q 0.08fF
C7775 BU_3VX2_71|A raven_soc_0|ext_clk 0.01fF
C7776 IN_3VX2_1|A raven_soc_0|gpio_in<7> 0.01fF
C7777 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<9> 2.39fF
C7778 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<14> 0.39fF
C7779 LS_3VX2_3|A raven_soc_0|flash_io3_di 0.01fF
C7780 BU_3VX2_0|Q raven_soc_0|flash_io1_do 0.03fF
C7781 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<11> 52.93fF
C7782 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<10> 2.61fF
C7783 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pullup<5> 0.02fF
C7784 raven_soc_0|gpio_outenb<15> raven_soc_0|ext_clk 0.01fF
C7785 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<12> 0.02fF
C7786 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<15> 0.02fF
C7787 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<20> 1.56fF
C7788 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<0> 0.02fF
C7789 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<28> 37.02fF
C7790 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<23> 4.36fF
C7791 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<19> 0.01fF
C7792 BU_3VX2_12|A BU_3VX2_26|A 0.01fF
C7793 LS_3VX2_12|A LS_3VX2_17|A 0.01fF
C7794 LS_3VX2_8|A BU_3VX2_62|Q 0.35fF
C7795 LOGIC0_3V_4|Q raven_soc_0|gpio_out<15> 25.54fF
C7796 BU_3VX2_13|A raven_soc_0|flash_io1_oeb 0.01fF
C7797 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pulldown<7> 0.02fF
C7798 BU_3VX2_33|A raven_soc_0|flash_io0_do 0.19fF
C7799 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<8> 0.14fF
C7800 VDD raven_padframe_0|BBCUD4F_8|GNDO 0.07fF
C7801 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<9> 4.56fF
C7802 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<14> 1.01fF
C7803 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_out<14> 0.47fF
C7804 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pullup<6> 0.02fF
C7805 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pulldown<6> 0.02fF
C7806 raven_soc_0|gpio_pulldown<9> BU_3VX2_71|Q 0.01fF
C7807 raven_soc_0|ram_wenb raven_soc_0|ram_addr<5> 0.01fF
C7808 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<17> 2.16fF
C7809 raven_soc_0|gpio_pulldown<8> vdd 0.31fF
C7810 raven_soc_0|gpio_pulldown<11> apllc03_1v8_0|CLK 0.20fF
C7811 raven_padframe_0|BBCUD4F_6|VDDR raven_padframe_0|BBCUD4F_6|GNDR 0.68fF
C7812 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<16> 6.15fF
C7813 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<18> 2.27fF
C7814 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<2> 3.53fF
C7815 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<12> 0.43fF
C7816 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<8> 13.39fF
C7817 BU_3VX2_68|Q BU_3VX2_65|Q 10.87fF
C7818 BU_3VX2_64|Q BU_3VX2_5|Q 0.90fF
C7819 raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<2> 44.15fF
C7820 BU_3VX2_73|Q BU_3VX2_57|Q 0.01fF
C7821 AMUX4_3V_3|SEL[0] BU_3VX2_33|Q 0.78fF
C7822 raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<8> 2.43fF
C7823 BU_3VX2_7|A BU_3VX2_21|A 0.41fF
C7824 raven_padframe_0|FILLER40F_0|GNDR raven_padframe_0|FILLER40F_0|VDDO 0.09fF
C7825 raven_padframe_0|CORNERESDF_2|GNDR raven_padframe_0|CORNERESDF_2|VDDO 0.09fF
C7826 LS_3VX2_8|A LS_3VX2_5|A 21.48fF
C7827 raven_padframe_0|APR00DF_1|VDDR adc_low 0.01fF
C7828 BU_3VX2_4|A BU_3VX2_27|A 0.01fF
C7829 BU_3VX2_63|A BU_3VX2_14|A 0.01fF
C7830 BU_3VX2_12|A BU_3VX2_11|A 36.80fF
C7831 raven_padframe_0|APR00DF_3|VDDO raven_padframe_0|APR00DF_3|GNDO 2.28fF
C7832 raven_padframe_0|FILLER02F_0|VDDO raven_padframe_0|FILLER02F_0|GNDO 2.32fF
C7833 LOGIC0_3V_4|Q raven_soc_0|gpio_in<5> 0.08fF
C7834 raven_soc_0|irq_pin LS_3VX2_15|A 0.01fF
C7835 raven_soc_0|ram_wdata<17> vdd 1.28fF
C7836 LS_3VX2_11|A LS_3VX2_11|Q 0.05fF
C7837 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<12> 0.01fF
C7838 BU_3VX2_67|A BU_3VX2_36|A 3.28fF
C7839 IN_3VX2_1|A raven_soc_0|gpio_out<7> 0.01fF
C7840 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<8> 0.01fF
C7841 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<7> 0.01fF
C7842 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_outenb<15> 1.05fF
C7843 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<14> 1.90fF
C7844 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<11> 4.57fF
C7845 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<6> 0.01fF
C7846 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<12> 26.18fF
C7847 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<13> 7.08fF
C7848 BU_3VX2_2|A BU_3VX2_35|Q 0.02fF
C7849 raven_soc_0|gpio_pullup<0> BU_3VX2_40|Q 0.02fF
C7850 raven_padframe_0|BBCUD4F_7|VDDR raven_padframe_0|BBCUD4F_7|GNDO 0.13fF
C7851 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io0_oeb 129.50fF
C7852 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<1> 4.34fF
C7853 BU_3VX2_21|Q BU_3VX2_32|Q 3.33fF
C7854 raven_soc_0|flash_io1_do raven_soc_0|flash_io3_di 76.54fF
C7855 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<17> 0.26fF
C7856 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<27> 0.06fF
C7857 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<31> 5.29fF
C7858 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<9> 0.87fF
C7859 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<24> 0.39fF
C7860 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<2> 93.51fF
C7861 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<10> 2.95fF
C7862 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<29> 0.06fF
C7863 BU_3VX2_2|Q BU_3VX2_11|Q 3.93fF
C7864 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<7> 0.64fF
C7865 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<22> 0.02fF
C7866 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<14> 0.03fF
C7867 raven_soc_0|flash_io3_do raven_soc_0|flash_io0_do 74.70fF
C7868 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<4> 87.06fF
C7869 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<23> 0.01fF
C7870 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<30> 6.10fF
C7871 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<2> 0.01fF
C7872 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<13> 4.56fF
C7873 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<25> 0.01fF
C7874 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<26> 0.01fF
C7875 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<21> 0.01fF
C7876 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<19> 0.01fF
C7877 BU_3VX2_11|Q BU_3VX2_10|Q 70.10fF
C7878 BU_3VX2_32|Q BU_3VX2_8|Q 0.67fF
C7879 BU_3VX2_4|Q BU_3VX2_22|Q 0.54fF
C7880 raven_soc_0|flash_io0_do AMUX4_3V_4|AIN3 1.27fF
C7881 BU_3VX2_60|Q vdd 1.95fF
C7882 BU_3VX2_29|Q BU_3VX2_27|Q 223.97fF
C7883 BU_3VX2_6|A raven_soc_0|flash_io0_oeb 0.01fF
C7884 BU_3VX2_38|A raven_soc_0|flash_io3_oeb 0.01fF
C7885 BU_3VX2_17|A VDD3V3 0.45fF
C7886 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<3> 0.94fF
C7887 IN_3VX2_1|A BU_3VX2_49|Q 5.70fF
C7888 LS_3VX2_4|A BU_3VX2_62|Q 0.31fF
C7889 BU_3VX2_28|A BU_3VX2_26|Q 0.03fF
C7890 raven_soc_0|gpio_pulldown<13> BU_3VX2_24|Q 0.01fF
C7891 BU_3VX2_71|Q raven_soc_0|flash_io0_di 12.40fF
C7892 raven_padframe_0|GNDORPADF_7|VDDR raven_padframe_0|GNDORPADF_7|VDDO 0.06fF
C7893 raven_soc_0|flash_clk BU_3VX2_11|Q 0.03fF
C7894 BU_3VX2_2|A BU_3VX2_38|A 10.23fF
C7895 LS_3VX2_5|A LS_3VX2_4|A 55.81fF
C7896 VDD raven_padframe_0|APR00DF_1|GNDO 0.07fF
C7897 LS_3VX2_6|A LS_3VX2_15|A 0.02fF
C7898 BU_3VX2_0|Q raven_soc_0|ram_rdata<31> 4.03fF
C7899 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<10> 0.01fF
C7900 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<11> 0.02fF
C7901 raven_soc_0|gpio_outenb<2> BU_3VX2_28|Q 0.01fF
C7902 raven_soc_0|gpio_pullup<1> BU_3VX2_24|Q 0.01fF
C7903 BU_3VX2_44|A LS_3VX2_27|Q 0.29fF
C7904 BU_3VX2_43|A LS_3VX2_21|Q 1.20fF
C7905 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<1> 127.86fF
C7906 LS_3VX2_14|A LS_3VX2_14|Q 0.05fF
C7907 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<9> 0.05fF
C7908 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_outenb<0> 9.54fF
C7909 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<5> 0.26fF
C7910 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<12> 0.01fF
C7911 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<8> 0.38fF
C7912 BU_3VX2_63|Q BU_3VX2_71|Q 87.46fF
C7913 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<8> 0.01fF
C7914 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<9> 20.02fF
C7915 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<14> 46.81fF
C7916 raven_padframe_0|FILLER10F_0|VDDR raven_padframe_0|FILLER10F_0|GNDO 0.13fF
C7917 raven_soc_0|flash_io1_do raven_soc_0|irq_pin 0.01fF
C7918 raven_soc_0|gpio_pulldown<7> VDD3V3 0.07fF
C7919 raven_soc_0|irq_pin AMUX4_3V_1|SEL[1] 0.01fF
C7920 BU_3VX2_73|Q LS_3VX2_16|A 0.01fF
C7921 BU_3VX2_65|Q BU_3VX2_24|Q 0.48fF
C7922 BU_3VX2_9|Q vdd 1.84fF
C7923 BU_3VX2_15|Q vdd 1.22fF
C7924 BU_3VX2_69|Q BU_3VX2_25|Q 0.33fF
C7925 BU_3VX2_64|Q BU_3VX2_28|Q 0.62fF
C7926 BU_3VX2_31|Q BU_3VX2_23|Q 3.50fF
C7927 BU_3VX2_35|Q apllc03_1v8_0|CLK 0.01fF
C7928 BU_3VX2_23|A BU_3VX2_3|A 0.01fF
C7929 BU_3VX2_23|A BU_3VX2_15|A 2.60fF
C7930 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<11> 2.05fF
C7931 BU_3VX2_72|A BU_3VX2_31|A 0.01fF
C7932 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<3> 0.99fF
C7933 BU_3VX2_12|A VDD3V3 0.46fF
C7934 raven_soc_0|ram_addr<9> raven_soc_0|ram_addr<0> 4.93fF
C7935 raven_soc_0|ram_wdata<22> raven_soc_0|ram_rdata<15> 2.41fF
C7936 raven_soc_0|ram_wdata<31> raven_soc_0|ram_rdata<13> 0.49fF
C7937 raven_soc_0|ram_wdata<29> raven_soc_0|ram_addr<0> 0.01fF
C7938 raven_soc_0|ram_wdata<25> raven_soc_0|ram_rdata<16> 0.01fF
C7939 raven_soc_0|flash_io0_oeb BU_3VX2_25|Q 0.01fF
C7940 BU_3VX2_53|Q LS_3VX2_27|A 0.05fF
C7941 BU_3VX2_51|A BU_3VX2_51|Q 0.10fF
C7942 BU_3VX2_55|A BU_3VX2_58|Q 0.02fF
C7943 raven_soc_0|flash_io2_oeb BU_3VX2_29|Q 0.01fF
C7944 BU_3VX2_60|A BU_3VX2_59|Q 0.03fF
C7945 raven_soc_0|flash_io3_oeb BU_3VX2_23|Q 0.01fF
C7946 raven_soc_0|flash_io2_do BU_3VX2_27|Q 0.01fF
C7947 raven_padframe_0|BT4FC_0|GNDR raven_padframe_0|BT4FC_0|GNDO 0.81fF
C7948 raven_padframe_0|ICF_0|GNDR raven_padframe_0|ICF_0|VDDO 0.09fF
C7949 raven_padframe_0|BBCUD4F_9|GNDR raven_padframe_0|BBCUD4F_9|GNDO 0.81fF
C7950 BU_3VX2_35|A raven_soc_0|flash_csb 0.01fF
C7951 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<6> 0.53fF
C7952 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<15> 0.01fF
C7953 BU_3VX2_24|A raven_soc_0|ext_clk 0.01fF
C7954 BU_3VX2_20|A BU_3VX2_20|Q 0.08fF
C7955 BU_3VX2_63|A raven_soc_0|flash_io1_do 0.01fF
C7956 VDD raven_padframe_0|BBCUD4F_13|GNDO 0.07fF
C7957 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<15> 17.41fF
C7958 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<5> 0.02fF
C7959 BU_3VX2_0|Q raven_soc_0|gpio_in<10> 0.09fF
C7960 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<14> 0.02fF
C7961 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<9> 35.38fF
C7962 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<12> 0.02fF
C7963 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<13> 0.02fF
C7964 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<28> 61.13fF
C7965 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<0> 1.76fF
C7966 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<19> 51.43fF
C7967 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<23> 0.02fF
C7968 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<20> 21.19fF
C7969 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<11> 0.01fF
C7970 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<3> 1.03fF
C7971 BU_3VX2_8|A raven_soc_0|flash_io0_do 0.01fF
C7972 LOGIC0_3V_4|Q raven_soc_0|gpio_in<6> 0.08fF
C7973 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<6> 0.83fF
C7974 LS_3VX2_6|A AMUX4_3V_1|SEL[1] 18.62fF
C7975 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<13> 0.01fF
C7976 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<14> 0.02fF
C7977 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pulldown<6> 0.02fF
C7978 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<5> 0.01fF
C7979 raven_spi_0|sdo_enb raven_soc_0|flash_io2_di 1.66fF
C7980 BU_3VX2_27|A raven_soc_0|flash_io0_oeb 6.70fF
C7981 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pulldown<7> 2.60fF
C7982 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<14> 0.02fF
C7983 BU_3VX2_33|A raven_soc_0|flash_io1_di 1.66fF
C7984 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<8> 9.07fF
C7985 raven_padframe_0|FILLER20F_3|VDDR raven_padframe_0|FILLER20F_3|GNDO 0.13fF
C7986 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<4> 19.26fF
C7987 LS_3VX2_7|A LS_3VX2_6|A 53.44fF
C7988 LOGIC0_3V_4|Q raven_soc_0|gpio_out<10> 0.01fF
C7989 raven_soc_0|gpio_out<2> BU_3VX2_71|Q 0.30fF
C7990 raven_soc_0|ram_wdata<18> vdd 0.63fF
C7991 raven_soc_0|ram_wdata<8> vdd 0.83fF
C7992 BU_3VX2_55|Q BU_3VX2_43|Q 0.02fF
C7993 BU_3VX2_54|A BU_3VX2_53|Q 0.03fF
C7994 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<5> 0.01fF
C7995 BU_3VX2_3|A IN_3VX2_1|A 0.01fF
C7996 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<0> 159.97fF
C7997 BU_3VX2_15|A IN_3VX2_1|A 0.01fF
C7998 raven_soc_0|gpio_outenb<3> BU_3VX2_63|Q 0.01fF
C7999 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<14> 0.06fF
C8000 IN_3VX2_1|A raven_soc_0|gpio_outenb<7> 0.01fF
C8001 raven_soc_0|gpio_in<0> BU_3VX2_0|Q 0.01fF
C8002 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<2> 12.30fF
C8003 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<11> 0.01fF
C8004 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<15> 0.05fF
C8005 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<14> 7.91fF
C8006 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<12> 38.04fF
C8007 BU_3VX2_0|Q raven_soc_0|flash_csb 0.01fF
C8008 raven_soc_0|gpio_out<1> BU_3VX2_27|Q 0.03fF
C8009 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<2> 8.80fF
C8010 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<4> 0.06fF
C8011 raven_soc_0|flash_io3_do raven_soc_0|flash_io1_di 75.51fF
C8012 BU_3VX2_66|Q BU_3VX2_14|Q 16.79fF
C8013 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<25> 0.14fF
C8014 raven_soc_0|flash_io2_do raven_soc_0|flash_io2_oeb 59.99fF
C8015 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<14> 0.02fF
C8016 BU_3VX2_15|Q BU_3VX2_70|Q 0.24fF
C8017 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<26> 0.73fF
C8018 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<6> 0.06fF
C8019 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<18> 1.13fF
C8020 BU_3VX2_19|Q BU_3VX2_32|Q 0.04fF
C8021 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<19> 3.48fF
C8022 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<8> 0.48fF
C8023 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<15> 12.54fF
C8024 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<2> 1.79fF
C8025 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<8> 0.07fF
C8026 BU_3VX2_13|Q BU_3VX2_37|Q 2.75fF
C8027 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<13> 0.01fF
C8028 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<4> 0.01fF
C8029 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<21> 3.96fF
C8030 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<6> 3.38fF
C8031 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<24> 4.03fF
C8032 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<2> 0.01fF
C8033 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<10> 0.01fF
C8034 BU_3VX2_3|Q BU_3VX2_22|Q 19.56fF
C8035 BU_3VX2_14|Q BU_3VX2_20|Q 5.88fF
C8036 BU_3VX2_36|Q BU_3VX2_68|Q 3.85fF
C8037 BU_3VX2_70|Q BU_3VX2_9|Q 2.86fF
C8038 BU_3VX2_23|Q apllc03_1v8_0|CLK 0.85fF
C8039 LS_3VX2_20|A BU_3VX2_47|Q 24.36fF
C8040 BU_3VX2_62|Q vdd 2.74fF
C8041 BU_3VX2_25|Q BU_3VX2_29|Q 64.62fF
C8042 BU_3VX2_44|Q BU_3VX2_45|Q 218.47fF
C8043 apllc03_1v8_0|B_VCO BU_3VX2_28|Q 0.39fF
C8044 BU_3VX2_26|Q apllc03_1v8_0|B_CP 1.29fF
C8045 raven_padframe_0|FILLER50F_1|VDDR raven_padframe_0|FILLER50F_1|VDDO 0.06fF
C8046 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<8> 0.01fF
C8047 LOGIC0_3V_4|Q raven_soc_0|gpio_in<3> 0.08fF
C8048 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_in<0> 137.27fF
C8049 raven_padframe_0|CORNERESDF_0|VDDO raven_padframe_0|CORNERESDF_0|GNDO 2.28fF
C8050 LOGIC0_3V_4|Q raven_soc_0|gpio_out<9> 0.01fF
C8051 raven_spi_0|SDO raven_soc_0|flash_io1_do 0.55fF
C8052 BU_3VX2_6|A raven_soc_0|flash_io2_do 0.02fF
C8053 BU_3VX2_73|A AMUX4_3V_4|AIN3 0.03fF
C8054 BU_3VX2_16|A raven_soc_0|ext_clk 0.13fF
C8055 raven_padframe_0|FILLER20F_1|VDDR raven_padframe_0|FILLER20F_1|GNDO 0.13fF
C8056 LS_3VX2_14|A BU_3VX2_51|Q 6.16fF
C8057 BU_3VX2_29|A raven_soc_0|ext_clk 0.01fF
C8058 LS_3VX2_5|A vdd 3.92fF
C8059 BU_3VX2_36|A BU_3VX2_33|Q 0.03fF
C8060 raven_soc_0|gpio_out<4> apllc03_1v8_0|CLK 0.01fF
C8061 LS_3VX2_3|A BU_3VX2_26|Q 0.01fF
C8062 raven_padframe_0|BBCUD4F_5|VDDR raven_padframe_0|BBCUD4F_5|GNDR 0.68fF
C8063 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<17> 44.54fF
C8064 BU_3VX2_22|A BU_3VX2_22|Q 0.08fF
C8065 LS_3VX2_9|A LS_3VX2_19|A 0.01fF
C8066 BU_3VX2_37|A raven_soc_0|ext_clk 0.01fF
C8067 LS_3VX2_9|A BU_3VX2_52|Q 26.24fF
C8068 AMUX4_3V_0|AIN1 AMUX4_3V_4|AIN2 1.09fF
C8069 BU_3VX2_4|A BU_3VX2_37|Q 0.02fF
C8070 LS_3VX2_12|A BU_3VX2_42|Q 5.60fF
C8071 BU_3VX2_11|A BU_3VX2_10|Q 0.16fF
C8072 BU_3VX2_26|A raven_soc_0|flash_clk 4.68fF
C8073 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<15> 0.02fF
C8074 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<13> 10.40fF
C8075 BU_3VX2_0|Q raven_soc_0|ram_rdata<30> 3.63fF
C8076 raven_soc_0|gpio_outenb<2> vdd 0.24fF
C8077 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_0|PO 0.04fF
C8078 VDD raven_padframe_0|APR00DF_0|VDDR 0.71fF
C8079 BU_3VX2_9|A BU_3VX2_26|A 0.01fF
C8080 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<10> 0.05fF
C8081 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<9> 0.46fF
C8082 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<7> 0.24fF
C8083 BU_3VX2_11|A raven_soc_0|flash_clk 0.01fF
C8084 raven_soc_0|gpio_in<0> raven_soc_0|flash_io3_di 0.22fF
C8085 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<6> 0.01fF
C8086 raven_soc_0|gpio_in<3> raven_soc_0|flash_io1_oeb 0.01fF
C8087 BU_3VX2_14|A BU_3VX2_11|Q 0.02fF
C8088 BU_3VX2_63|Q raven_soc_0|gpio_pullup<14> 0.01fF
C8089 raven_soc_0|flash_csb raven_soc_0|flash_io3_di 13.50fF
C8090 raven_soc_0|gpio_in<10> raven_soc_0|irq_pin 0.01fF
C8091 AMUX4_3V_0|SEL[1] BU_3VX2_56|Q 0.43fF
C8092 BU_3VX2_64|Q vdd 2.67fF
C8093 LS_3VX2_11|A LS_3VX2_8|A 33.62fF
C8094 LS_3VX2_13|Q LS_3VX2_9|Q 0.55fF
C8095 BU_3VX2_9|A BU_3VX2_11|A 7.68fF
C8096 BU_3VX2_0|A BU_3VX2_33|A 1.86fF
C8097 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<2> 4.14fF
C8098 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<5> 2.32fF
C8099 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<2> 105.76fF
C8100 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<16> 0.18fF
C8101 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<0> 19.92fF
C8102 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<15> 5.87fF
C8103 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<16> 6.67fF
C8104 raven_soc_0|ram_wdata<19> raven_soc_0|ram_rdata<13> 0.04fF
C8105 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<29> 0.01fF
C8106 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<31> 0.01fF
C8107 BU_3VX2_48|A LS_3VX2_27|Q 0.12fF
C8108 BU_3VX2_49|A BU_3VX2_42|A 0.15fF
C8109 BU_3VX2_47|A LS_3VX2_20|Q 0.22fF
C8110 BU_3VX2_41|A BU_3VX2_44|A 1.06fF
C8111 BU_3VX2_62|A BU_3VX2_62|Q 0.10fF
C8112 BU_3VX2_48|A BU_3VX2_48|Q 0.10fF
C8113 BU_3VX2_51|A BU_3VX2_49|Q 0.04fF
C8114 BU_3VX2_60|A BU_3VX2_61|Q 0.14fF
C8115 raven_soc_0|flash_io3_do BU_3VX2_28|Q 0.01fF
C8116 raven_soc_0|flash_io1_do BU_3VX2_26|Q 0.01fF
C8117 raven_soc_0|flash_io2_do BU_3VX2_25|Q 0.01fF
C8118 BU_3VX2_45|Q vdd 1.78fF
C8119 BU_3VX2_3|A BU_3VX2_25|A 0.01fF
C8120 BU_3VX2_25|A BU_3VX2_15|A 2.05fF
C8121 LS_3VX2_11|Q LS_3VX2_10|Q 3.65fF
C8122 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<14> 0.01fF
C8123 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<11> 0.48fF
C8124 raven_padframe_0|axtoc02_3v3_0|m4_0_28769# raven_padframe_0|axtoc02_3v3_0|m4_0_22024# 0.06fF
C8125 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<12> 7.42fF
C8126 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<13> 13.37fF
C8127 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<14> 0.02fF
C8128 BU_3VX2_10|A raven_soc_0|flash_io3_do 0.03fF
C8129 BU_3VX2_8|A BU_3VX2_5|Q 0.02fF
C8130 IN_3VX2_1|Q raven_soc_0|irq_pin 159.68fF
C8131 LS_3VX2_10|A BU_3VX2_55|Q 9.53fF
C8132 LS_3VX2_3|Q raven_soc_0|ext_clk 0.01fF
C8133 BU_3VX2_31|A BU_3VX2_31|Q 0.08fF
C8134 raven_padframe_0|POWERCUTVDD3FC_0|VDDR raven_padframe_0|POWERCUTVDD3FC_0|GNDR 0.64fF
C8135 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<5> 0.01fF
C8136 raven_soc_0|gpio_pullup<3> BU_3VX2_40|Q 0.33fF
C8137 BU_3VX2_0|Q raven_soc_0|gpio_in<13> 0.35fF
C8138 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<7> 0.55fF
C8139 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<6> 0.01fF
C8140 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<9> 99.03fF
C8141 raven_soc_0|gpio_pullup<4> VDD3V3 0.09fF
C8142 raven_padframe_0|FILLER02F_1|VDDR raven_padframe_0|FILLER02F_1|VDDO 0.06fF
C8143 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<28> 0.01fF
C8144 BU_3VX2_71|Q BU_3VX2_24|Q 1.86fF
C8145 raven_soc_0|gpio_out<14> BU_3VX2_28|Q 0.01fF
C8146 BU_3VX2_32|Q BU_3VX2_27|Q 0.13fF
C8147 BU_3VX2_36|Q BU_3VX2_24|Q 1.33fF
C8148 BU_3VX2_4|Q apllc03_1v8_0|CLK 0.01fF
C8149 BU_3VX2_32|A BU_3VX2_32|Q 0.08fF
C8150 BU_3VX2_21|A BU_3VX2_22|Q 0.03fF
C8151 BU_3VX2_8|A raven_soc_0|flash_io1_di 0.01fF
C8152 BU_3VX2_20|A raven_soc_0|flash_io3_di 0.01fF
C8153 BU_3VX2_0|A raven_soc_0|flash_io3_do 7.81fF
C8154 BU_3VX2_18|A raven_soc_0|flash_io2_di 0.01fF
C8155 BU_3VX2_67|A VDD3V3 0.02fF
C8156 raven_padframe_0|BBC4F_3|VDDR raven_padframe_0|BBC4F_3|GNDO 0.13fF
C8157 LOGIC0_3V_4|Q raven_soc_0|ext_clk 0.08fF
C8158 VDD raven_padframe_0|ICF_0|GNDO 0.07fF
C8159 raven_soc_0|gpio_in<0> raven_soc_0|irq_pin 0.01fF
C8160 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<8> 0.06fF
C8161 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<10> 0.01fF
C8162 BU_3VX2_31|A raven_soc_0|flash_io3_oeb 20.06fF
C8163 LS_3VX2_3|A raven_soc_0|gpio_outenb<13> 0.32fF
C8164 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<6> 0.10fF
C8165 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<14> 15.39fF
C8166 BU_3VX2_27|A raven_soc_0|flash_io2_do 3.40fF
C8167 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pulldown<7> 7.37fF
C8168 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<12> 0.31fF
C8169 BU_3VX2_0|Q BU_3VX2_14|Q 0.01fF
C8170 BU_3VX2_2|A BU_3VX2_31|A 0.01fF
C8171 LS_3VX2_11|A LS_3VX2_4|A 18.23fF
C8172 BU_3VX2_28|A BU_3VX2_26|A 20.18fF
C8173 LS_3VX2_9|A BU_3VX2_58|Q 8.66fF
C8174 LS_3VX2_8|A LS_3VX2_21|A 7.31fF
C8175 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<9> 0.35fF
C8176 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<14> 0.01fF
C8177 raven_soc_0|gpio_out<11> BU_3VX2_27|Q 0.01fF
C8178 raven_padframe_0|FILLER20F_0|VDDR VDD 0.71fF
C8179 BU_3VX2_56|A BU_3VX2_55|Q 0.03fF
C8180 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<7> 0.01fF
C8181 BU_3VX2_19|A BU_3VX2_17|A 12.42fF
C8182 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<10> 0.01fF
C8183 BU_3VX2_63|A raven_soc_0|flash_csb 0.01fF
C8184 BU_3VX2_28|A BU_3VX2_11|A 0.01fF
C8185 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<15> 0.01fF
C8186 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<3> 0.01fF
C8187 IN_3VX2_1|A raven_soc_0|gpio_pullup<9> 0.01fF
C8188 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<9> 0.01fF
C8189 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<15> 1.20fF
C8190 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<5> 0.47fF
C8191 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_outenb<6> 0.03fF
C8192 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<12> 0.11fF
C8193 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<12> 11.34fF
C8194 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<7> 1.22fF
C8195 raven_soc_0|gpio_out<1> BU_3VX2_25|Q 0.01fF
C8196 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<22> 23.97fF
C8197 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<23> 10.77fF
C8198 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<5> 4.34fF
C8199 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<20> 3.66fF
C8200 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<8> 0.02fF
C8201 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<9> 0.05fF
C8202 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<24> 0.22fF
C8203 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<10> 1.01fF
C8204 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<18> 0.25fF
C8205 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<13> 0.01fF
C8206 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<14> 13.52fF
C8207 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<0> 0.07fF
C8208 BU_3VX2_16|Q BU_3VX2_14|Q 22.82fF
C8209 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<25> 4.45fF
C8210 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<15> 1.58fF
C8211 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<2> 0.01fF
C8212 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<12> 0.10fF
C8213 raven_soc_0|ext_clk raven_soc_0|flash_io1_oeb 27.03fF
C8214 BU_3VX2_14|Q BU_3VX2_30|Q 0.14fF
C8215 BU_3VX2_70|Q BU_3VX2_64|Q 3.44fF
C8216 BU_3VX2_37|Q BU_3VX2_69|Q 0.11fF
C8217 AMUX4_3V_4|AIN3 comp_inp 183.79fF
C8218 raven_padframe_0|FILLER20F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C8219 raven_soc_0|flash_clk VDD3V3 12.90fF
C8220 BU_3VX2_42|Q BU_3VX2_46|Q 19.29fF
C8221 LOGIC0_3V_0|Q BU_3VX2_33|A 1.93fF
C8222 LOGIC0_3V_1|Q LOGIC0_3V_2|Q 20.99fF
C8223 vdd apllc03_1v8_0|B_VCO 5.17fF
C8224 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<10> 0.01fF
C8225 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<1> 2.07fF
C8226 AMUX4_3V_1|AIN1 BU_3VX2_61|A 0.02fF
C8227 BU_3VX2_9|A VDD3V3 0.14fF
C8228 VDD raven_padframe_0|BT4F_1|GNDR 0.16fF
C8229 LS_3VX2_14|A BU_3VX2_49|Q 5.11fF
C8230 VDD raven_padframe_0|BBCUD4F_1|GNDR 0.16fF
C8231 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<1> 0.44fF
C8232 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<27> 0.02fF
C8233 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<22> 0.02fF
C8234 BU_3VX2_71|Q raven_soc_0|gpio_out<15> 0.09fF
C8235 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<31> 3.45fF
C8236 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<19> 0.01fF
C8237 raven_soc_0|ram_rdata<23> raven_soc_0|ram_wdata<25> 0.01fF
C8238 LS_3VX2_9|A LS_3VX2_22|A 8.00fF
C8239 BU_3VX2_2|A BU_3VX2_3|Q 0.03fF
C8240 BU_3VX2_15|A BU_3VX2_13|Q 0.03fF
C8241 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<14> 0.02fF
C8242 BU_3VX2_63|Q raven_soc_0|gpio_in<9> 0.01fF
C8243 BU_3VX2_31|A apllc03_1v8_0|CLK 4.14fF
C8244 raven_soc_0|gpio_pulldown<1> BU_3VX2_28|Q 0.01fF
C8245 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<5> 0.01fF
C8246 AMUX2_3V_0|SEL VDD3V3 0.74fF
C8247 BU_3VX2_33|A vdd 0.06fF
C8248 raven_soc_0|gpio_in<5> BU_3VX2_71|Q 0.28fF
C8249 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<10> 0.67fF
C8250 raven_padframe_0|ICFC_1|GNDR raven_padframe_0|ICFC_1|GNDO 0.81fF
C8251 BU_3VX2_10|A BU_3VX2_8|A 10.86fF
C8252 BU_3VX2_20|A BU_3VX2_63|A 0.01fF
C8253 BU_3VX2_19|A BU_3VX2_12|A 2.44fF
C8254 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<12> 0.35fF
C8255 raven_soc_0|gpio_outenb<1> BU_3VX2_0|Q 0.30fF
C8256 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<9> 0.01fF
C8257 BU_3VX2_22|A raven_soc_0|flash_io3_oeb 0.01fF
C8258 BU_3VX2_71|A raven_soc_0|flash_io2_di 0.01fF
C8259 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<8> 0.36fF
C8260 raven_padframe_0|BBCUD4F_15|VDDR raven_padframe_0|BBCUD4F_15|GNDR 0.68fF
C8261 LOGIC0_3V_4|Q raven_padframe_0|BBC4F_3|PO 0.04fF
C8262 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<3> 0.15fF
C8263 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<6> 0.01fF
C8264 LS_3VX2_18|Q acmpc01_3v3_0|IBN 4.15fF
C8265 raven_soc_0|gpio_in<13> raven_soc_0|irq_pin 0.01fF
C8266 BU_3VX2_56|Q BU_3VX2_49|Q 0.03fF
C8267 BU_3VX2_3|A BU_3VX2_4|A 20.73fF
C8268 BU_3VX2_8|A BU_3VX2_0|A 0.01fF
C8269 BU_3VX2_4|A BU_3VX2_15|A 0.93fF
C8270 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_outenb<1> 27.64fF
C8271 BU_3VX2_26|A BU_3VX2_14|A 1.67fF
C8272 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<7> 30.04fF
C8273 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<9> 2.84fF
C8274 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<31> 8.29fF
C8275 raven_soc_0|ram_rdata<25> raven_soc_0|ram_addr<0> 7.56fF
C8276 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<13> 0.28fF
C8277 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<29> 0.71fF
C8278 raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<25> 27.56fF
C8279 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<27> 7.46fF
C8280 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<19> 0.01fF
C8281 raven_soc_0|flash_io3_do vdd 2.57fF
C8282 raven_soc_0|gpio_in<12> BU_3VX2_27|Q 0.01fF
C8283 raven_soc_0|ser_tx BU_3VX2_55|Q 5.53fF
C8284 VDD3V3 BU_3VX2_61|Q 0.04fF
C8285 raven_soc_0|gpio_in<15> BU_3VX2_23|Q 0.01fF
C8286 raven_soc_0|gpio_in<10> BU_3VX2_26|Q 0.01fF
C8287 AMUX4_3V_4|AIN3 vdd 7.78fF
C8288 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<15> 0.01fF
C8289 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<2> 20.08fF
C8290 BU_3VX2_11|A BU_3VX2_14|A 6.87fF
C8291 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<12> 8.38fF
C8292 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<15> 0.02fF
C8293 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<11> 0.01fF
C8294 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<15> 0.02fF
C8295 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<5> 0.01fF
C8296 LS_3VX2_10|A BU_3VX2_57|Q 7.68fF
C8297 BU_3VX2_28|A VDD3V3 1.23fF
C8298 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<15> 0.67fF
C8299 LS_3VX2_24|A BU_3VX2_55|Q 0.02fF
C8300 raven_soc_0|gpio_pulldown<13> raven_soc_0|ext_clk 0.01fF
C8301 raven_soc_0|gpio_pulldown<5> BU_3VX2_40|Q 0.26fF
C8302 LS_3VX2_3|A raven_soc_0|gpio_in<8> 0.01fF
C8303 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<5> 0.01fF
C8304 raven_soc_0|gpio_out<14> vdd 0.17fF
C8305 raven_soc_0|gpio_pullup<14> BU_3VX2_24|Q 0.01fF
C8306 raven_soc_0|gpio_out<8> apllc03_1v8_0|CLK 0.01fF
C8307 LS_3VX2_21|A BU_3VX2_44|Q 8.16fF
C8308 BU_3VX2_37|Q BU_3VX2_29|Q 0.01fF
C8309 BU_3VX2_3|Q apllc03_1v8_0|CLK 0.01fF
C8310 BU_3VX2_40|A raven_soc_0|flash_io3_do 0.01fF
C8311 LS_3VX2_11|A vdd 2.57fF
C8312 raven_padframe_0|BT4F_1|VDDR raven_padframe_0|BT4F_1|GNDR 0.68fF
C8313 BU_3VX2_17|A BU_3VX2_18|Q 0.03fF
C8314 raven_soc_0|gpio_in<2> raven_soc_0|flash_io3_do 8.19fF
C8315 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<9> 0.22fF
C8316 BU_3VX2_0|Q raven_soc_0|gpio_pulldown<3> 0.17fF
C8317 raven_soc_0|gpio_pullup<1> raven_soc_0|ext_clk 0.03fF
C8318 LS_3VX2_3|A raven_soc_0|gpio_pullup<13> 0.17fF
C8319 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<0> 0.18fF
C8320 BU_3VX2_50|A BU_3VX2_45|A 0.59fF
C8321 BU_3VX2_48|A BU_3VX2_41|A 3.29fF
C8322 BU_3VX2_46|A adc0_data<5> 0.03fF
C8323 BU_3VX2_50|A BU_3VX2_47|Q 0.02fF
C8324 raven_padframe_0|BBCUD4F_11|VDDO raven_padframe_0|BBCUD4F_11|GNDO 2.28fF
C8325 BU_3VX2_23|A raven_soc_0|flash_io0_di 0.01fF
C8326 LS_3VX2_9|A BU_3VX2_60|Q 7.09fF
C8327 BU_3VX2_21|A raven_soc_0|flash_io3_oeb 0.01fF
C8328 LS_3VX2_9|Q LS_3VX2_19|A 0.01fF
C8329 raven_soc_0|gpio_out<0> BU_3VX2_28|Q 0.01fF
C8330 BU_3VX2_31|A raven_soc_0|gpio_outenb<8> 0.01fF
C8331 raven_padframe_0|ICFC_1|VDDR raven_padframe_0|ICFC_1|GNDR 0.68fF
C8332 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<3> 0.99fF
C8333 VDD raven_padframe_0|APR00DF_6|GNDO 0.07fF
C8334 raven_padframe_0|ICF_0|VDDR raven_padframe_0|ICF_0|GNDR 0.68fF
C8335 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<14> 0.10fF
C8336 LS_3VX2_8|A LS_3VX2_27|A 8.48fF
C8337 raven_soc_0|gpio_in<0> BU_3VX2_26|Q 0.01fF
C8338 raven_soc_0|gpio_out<11> BU_3VX2_25|Q 0.01fF
C8339 raven_soc_0|gpio_out<12> BU_3VX2_28|Q 0.01fF
C8340 raven_soc_0|gpio_out<6> apllc03_1v8_0|CLK 0.01fF
C8341 raven_soc_0|gpio_out<13> BU_3VX2_23|Q 0.01fF
C8342 raven_soc_0|flash_csb BU_3VX2_26|Q 10.11fF
C8343 BU_3VX2_56|A BU_3VX2_57|Q 0.15fF
C8344 raven_soc_0|gpio_in<1> BU_3VX2_0|Q 0.01fF
C8345 VDD raven_padframe_0|BBCUD4F_10|VDDR 0.71fF
C8346 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<12> 0.01fF
C8347 LS_3VX2_12|Q LS_3VX2_13|A 0.16fF
C8348 IN_3VX2_1|A raven_soc_0|gpio_pulldown<9> 0.01fF
C8349 LS_3VX2_23|Q LS_3VX2_23|A 0.04fF
C8350 raven_soc_0|gpio_out<4> raven_soc_0|gpio_out<13> 3.49fF
C8351 raven_soc_0|gpio_pullup<0> BU_3VX2_63|Q 0.01fF
C8352 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<2> 0.69fF
C8353 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<9> 0.94fF
C8354 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<8> 0.53fF
C8355 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<12> 0.89fF
C8356 LS_3VX2_3|A raven_soc_0|gpio_out<5> 0.01fF
C8357 BU_3VX2_0|Q raven_soc_0|gpio_outenb<5> 0.01fF
C8358 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<10> 0.01fF
C8359 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<12> 10.27fF
C8360 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<7> 1.47fF
C8361 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<12> 36.42fF
C8362 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<9> 0.04fF
C8363 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<7> 8.21fF
C8364 AMUX4_3V_3|SEL[1] BU_3VX2_6|Q 0.20fF
C8365 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<10> 84.41fF
C8366 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<14> 0.03fF
C8367 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<12> 3.68fF
C8368 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<0> 0.67fF
C8369 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<1> 0.01fF
C8370 AMUX4_3V_3|SEL[1] BU_3VX2_7|Q 0.69fF
C8371 BU_3VX2_40|Q raven_soc_0|flash_io0_oeb 0.01fF
C8372 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<0> 18.79fF
C8373 raven_padframe_0|ICF_1|GNDR raven_padframe_0|ICF_1|VDDO 0.09fF
C8374 raven_padframe_0|FILLER20F_8|VDDO raven_padframe_0|FILLER20F_8|GNDO 2.28fF
C8375 raven_padframe_0|BBCUD4F_10|VDDR LOGIC0_3V_4|Q 0.01fF
C8376 LOGIC1_3V_0|Q LOGIC0_3V_3|Q 0.17fF
C8377 LS_3VX2_9|Q adc_low 0.12fF
C8378 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<10> 0.01fF
C8379 raven_padframe_0|aregc01_3v3_0|m4_92500_29057# raven_padframe_0|aregc01_3v3_0|m4_92500_22024# 0.02fF
C8380 raven_padframe_0|aregc01_3v3_0|m4_0_29057# raven_padframe_0|aregc01_3v3_0|VDDO 0.04fF
C8381 raven_padframe_0|aregc01_3v3_0|m4_0_29333# raven_padframe_0|aregc01_3v3_0|GNDO 0.12fF
C8382 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<14> 1.10fF
C8383 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<11> 7.69fF
C8384 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<19> 9.86fF
C8385 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<11> 0.47fF
C8386 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<23> 33.00fF
C8387 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<20> 7.01fF
C8388 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<10> 0.02fF
C8389 BU_3VX2_71|Q raven_soc_0|gpio_in<6> 0.02fF
C8390 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<28> 4.82fF
C8391 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_out<15> 230.48fF
C8392 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<26> 0.02fF
C8393 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<17> 0.01fF
C8394 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<19> 0.01fF
C8395 raven_soc_0|ram_rdata<9> vdd 0.21fF
C8396 raven_soc_0|ram_rdata<18> apllc03_1v8_0|CLK 0.01fF
C8397 LS_3VX2_21|A vdd 3.48fF
C8398 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<8> 0.01fF
C8399 BU_3VX2_8|A vdd 0.12fF
C8400 LS_3VX2_10|A LS_3VX2_16|A 0.01fF
C8401 BU_3VX2_65|A BU_3VX2_65|Q 0.08fF
C8402 BU_3VX2_26|A raven_soc_0|flash_io1_do 2.45fF
C8403 BU_3VX2_14|A VDD3V3 0.42fF
C8404 raven_soc_0|gpio_pulldown<1> vdd 0.21fF
C8405 raven_soc_0|gpio_pulldown<2> apllc03_1v8_0|CLK 0.01fF
C8406 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<31> 14.82fF
C8407 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<6> 22.97fF
C8408 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<10> 1.79fF
C8409 raven_soc_0|gpio_out<8> raven_soc_0|gpio_outenb<8> 73.59fF
C8410 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_out<14> 0.27fF
C8411 raven_soc_0|gpio_out<10> BU_3VX2_71|Q 0.66fF
C8412 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<5> 0.01fF
C8413 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<24> 0.01fF
C8414 raven_padframe_0|ICF_2|VDDO raven_padframe_0|ICF_2|GNDO 2.28fF
C8415 raven_padframe_0|BBCUD4F_14|GNDR raven_padframe_0|BBCUD4F_14|VDDO 0.09fF
C8416 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<4> 0.01fF
C8417 markings_0|efabless_logo_0|m1_3300_n1350# markings_0|efabless_logo_0|m1_6600_n2850# 0.35fF
C8418 raven_soc_0|gpio_in<1> raven_soc_0|flash_io3_di 0.28fF
C8419 BU_3VX2_24|A raven_soc_0|flash_io2_di 0.01fF
C8420 AMUX4_3V_3|AOUT raven_soc_0|flash_io2_oeb 0.74fF
C8421 BU_3VX2_3|A raven_soc_0|flash_io0_oeb 0.01fF
C8422 BU_3VX2_15|A raven_soc_0|flash_io0_oeb 0.01fF
C8423 IN_3VX2_1|A raven_soc_0|flash_io0_di 0.01fF
C8424 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<6> 0.47fF
C8425 BU_3VX2_11|A raven_soc_0|flash_io1_do 0.01fF
C8426 IN_3VX2_1|A BU_3VX2_46|Q 8.42fF
C8427 raven_soc_0|irq_pin LS_3VX2_20|A 0.01fF
C8428 VDD raven_padframe_0|BBCUD4F_4|VDDR 0.71fF
C8429 BU_3VX2_38|A BU_3VX2_71|A 0.01fF
C8430 BU_3VX2_8|A BU_3VX2_40|A 0.58fF
C8431 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_in<2> 15.25fF
C8432 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_out<2> 10.45fF
C8433 AMUX4_3V_0|AIN1 BU_3VX2_46|A 0.02fF
C8434 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<13> 0.01fF
C8435 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<7> 0.11fF
C8436 raven_soc_0|gpio_in<3> BU_3VX2_71|Q 0.18fF
C8437 raven_soc_0|gpio_out<6> raven_soc_0|gpio_outenb<8> 1.28fF
C8438 raven_soc_0|gpio_out<9> BU_3VX2_71|Q 0.01fF
C8439 BU_3VX2_2|Q BU_3VX2_21|Q 0.50fF
C8440 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<7> 0.01fF
C8441 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<17> 0.01fF
C8442 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<27> 8.73fF
C8443 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<25> 2.14fF
C8444 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<25> 0.01fF
C8445 raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<31> 0.01fF
C8446 BU_3VX2_13|Q BU_3VX2_17|Q 10.81fF
C8447 BU_3VX2_66|Q BU_3VX2_20|Q 0.01fF
C8448 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<13> 80.75fF
C8449 BU_3VX2_21|Q BU_3VX2_10|Q 2.98fF
C8450 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<26> 12.39fF
C8451 BU_3VX2_2|Q BU_3VX2_8|Q 8.66fF
C8452 BU_3VX2_10|Q BU_3VX2_8|Q 29.31fF
C8453 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<19> 0.29fF
C8454 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<21> 6.75fF
C8455 raven_soc_0|ram_wdata<1> raven_soc_0|ram_rdata<17> 0.13fF
C8456 BU_3VX2_73|Q BU_3VX2_52|Q 0.01fF
C8457 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<22> 8.17fF
C8458 raven_soc_0|ser_tx BU_3VX2_57|Q 6.71fF
C8459 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<25> 4.87fF
C8460 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<29> 0.01fF
C8461 LS_3VX2_15|Q LS_3VX2_17|A 0.01fF
C8462 raven_soc_0|ext_clk BU_3VX2_72|Q 0.69fF
C8463 VDD3V3 LS_3VX2_15|A 0.43fF
C8464 raven_soc_0|gpio_in<9> BU_3VX2_24|Q 0.01fF
C8465 raven_soc_0|gpio_in<14> BU_3VX2_23|Q 0.01fF
C8466 raven_soc_0|gpio_in<12> BU_3VX2_25|Q 0.01fF
C8467 raven_soc_0|gpio_in<13> BU_3VX2_26|Q 0.01fF
C8468 BU_3VX2_40|Q BU_3VX2_29|Q 2.37fF
C8469 LS_3VX2_17|Q vdd 0.04fF
C8470 BU_3VX2_23|A BU_3VX2_5|A 0.01fF
C8471 raven_padframe_0|BBCUD4F_4|VDDR LOGIC0_3V_4|Q 0.01fF
C8472 raven_padframe_0|APR00DF_2|GNDR raven_padframe_0|APR00DF_2|GNDO 0.81fF
C8473 raven_padframe_0|axtoc02_3v3_0|m4_0_29333# raven_padframe_0|axtoc02_3v3_0|m4_0_29057# 0.22fF
C8474 raven_padframe_0|axtoc02_3v3_0|m4_0_30133# raven_padframe_0|axtoc02_3v3_0|m4_0_28769# 0.02fF
C8475 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<7> 0.01fF
C8476 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<12> 12.63fF
C8477 LS_3VX2_24|A BU_3VX2_57|Q 0.02fF
C8478 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<14> 0.01fF
C8479 LS_3VX2_3|A VDD3V3 0.74fF
C8480 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<5> 0.01fF
C8481 BU_3VX2_1|Q raven_soc_0|flash_io1_di 0.01fF
C8482 BU_3VX2_14|Q BU_3VX2_26|Q 3.51fF
C8483 raven_soc_0|gpio_pulldown<6> apllc03_1v8_0|CLK 0.07fF
C8484 LS_3VX2_27|A BU_3VX2_44|Q 7.73fF
C8485 raven_soc_0|gpio_in<1> raven_soc_0|irq_pin 0.01fF
C8486 LOGIC1_3V_0|Q VDD3V3 0.06fF
C8487 BU_3VX2_9|A BU_3VX2_8|Q 0.16fF
C8488 IN_3VX2_1|Q AMUX4_3V_0|SEL[0] 6.71fF
C8489 VDD raven_padframe_0|FILLER50F_2|GNDO 0.07fF
C8490 VDD raven_padframe_0|FILLER20F_7|GNDO 0.07fF
C8491 adc_low BU_3VX2_73|Q 0.05fF
C8492 BU_3VX2_31|A raven_soc_0|gpio_in<15> 0.01fF
C8493 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<6> 0.01fF
C8494 raven_padframe_0|BBCUD4F_10|VDDR raven_padframe_0|BBCUD4F_10|GNDR 0.68fF
C8495 BU_3VX2_51|A BU_3VX2_49|A 4.42fF
C8496 raven_padframe_0|FILLER20F_0|GNDR raven_padframe_0|FILLER20F_0|GNDO 0.81fF
C8497 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<7> 0.15fF
C8498 LS_3VX2_9|A BU_3VX2_62|Q 3.05fF
C8499 BU_3VX2_19|A raven_soc_0|flash_clk 0.01fF
C8500 raven_soc_0|gpio_out<0> vdd 1.59fF
C8501 BU_3VX2_16|A raven_soc_0|flash_io2_di 0.08fF
C8502 LS_3VX2_9|Q LS_3VX2_22|A 0.01fF
C8503 LS_3VX2_12|A BU_3VX2_54|Q 6.82fF
C8504 BU_3VX2_17|A raven_soc_0|flash_io2_oeb 0.01fF
C8505 VDD raven_padframe_0|APR00DF_6|VDDR 0.71fF
C8506 raven_padframe_0|ICFC_2|VDDR raven_padframe_0|ICFC_2|GNDO 0.13fF
C8507 raven_padframe_0|ICFC_2|VDD3 raven_padframe_0|ICFC_2|GNDR 0.16fF
C8508 raven_padframe_0|POWERCUTVDD3FC_1|VDDR raven_padframe_0|POWERCUTVDD3FC_1|VDDO 0.06fF
C8509 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<10> 0.01fF
C8510 BU_3VX2_29|A raven_soc_0|flash_io2_di 0.01fF
C8511 raven_soc_0|gpio_out<12> vdd 0.18fF
C8512 VDD raven_padframe_0|FILLER10F_0|GNDO 0.07fF
C8513 raven_soc_0|gpio_outenb<12> BU_3VX2_28|Q 0.01fF
C8514 raven_soc_0|gpio_outenb<11> apllc03_1v8_0|CLK 0.01fF
C8515 raven_soc_0|gpio_outenb<15> BU_3VX2_23|Q 0.01fF
C8516 BU_3VX2_9|A BU_3VX2_19|A 1.22fF
C8517 BU_3VX2_6|A BU_3VX2_17|A 1.00fF
C8518 LS_3VX2_9|A LS_3VX2_5|A 157.25fF
C8519 IN_3VX2_1|Q analog_out 1.95fF
C8520 raven_soc_0|gpio_out<4> raven_soc_0|gpio_outenb<15> 1.13fF
C8521 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<3> 0.04fF
C8522 LS_3VX2_3|A raven_soc_0|gpio_outenb<6> 0.01fF
C8523 BU_3VX2_0|Q raven_soc_0|gpio_pullup<7> 0.01fF
C8524 BU_3VX2_37|A raven_soc_0|flash_io2_di 0.01fF
C8525 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<12> 7.64fF
C8526 BU_3VX2_25|A raven_soc_0|flash_io0_di 0.01fF
C8527 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<9> 0.02fF
C8528 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<10> 0.01fF
C8529 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<12> 62.21fF
C8530 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<8> 0.02fF
C8531 BU_3VX2_40|Q raven_soc_0|flash_io2_do 0.01fF
C8532 raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<10> 6.79fF
C8533 raven_soc_0|gpio_in<9> raven_soc_0|gpio_out<15> 0.01fF
C8534 raven_soc_0|flash_io1_do VDD3V3 11.87fF
C8535 LS_3VX2_17|Q BU_3VX2_62|A 2.81fF
C8536 VDD3V3 AMUX4_3V_1|SEL[1] 0.66fF
C8537 VDD raven_padframe_0|BT4F_0|VDDR 0.71fF
C8538 raven_padframe_0|BT4F_2|GNDR raven_padframe_0|BT4F_2|GNDO 0.81fF
C8539 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<2> 9.08fF
C8540 BU_3VX2_5|A IN_3VX2_1|A 0.01fF
C8541 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_in<3> 34.47fF
C8542 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<4> 0.01fF
C8543 IN_3VX2_1|A raven_soc_0|gpio_out<2> 0.01fF
C8544 BU_3VX2_31|A raven_soc_0|gpio_out<13> 0.01fF
C8545 raven_padframe_0|aregc01_3v3_0|m4_92500_31172# raven_padframe_0|aregc01_3v3_0|m4_92500_30653# 0.09fF
C8546 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<12> 0.04fF
C8547 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<7> 0.37fF
C8548 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<9> 0.02fF
C8549 BU_3VX2_69|A BU_3VX2_33|A 1.07fF
C8550 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<15> 0.76fF
C8551 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<10> 0.11fF
C8552 markings_0|efabless_logo_0|m1_6600_n9150# markings_0|efabless_logo_0|m1_4500_n11550# 0.31fF
C8553 BU_3VX2_68|A BU_3VX2_68|Q 0.08fF
C8554 LS_3VX2_7|A VDD3V3 0.52fF
C8555 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<9> 0.79fF
C8556 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<0> 0.12fF
C8557 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<20> 0.32fF
C8558 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<23> 0.14fF
C8559 BU_3VX2_71|Q raven_soc_0|ext_clk 20.28fF
C8560 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<6> 0.01fF
C8561 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<11> 3.17fF
C8562 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<13> 190.50fF
C8563 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<15> 0.02fF
C8564 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<10> 0.01fF
C8565 raven_soc_0|ser_tx LS_3VX2_16|A 26.68fF
C8566 BU_3VX2_73|Q BU_3VX2_58|Q 0.01fF
C8567 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<8> 0.01fF
C8568 raven_soc_0|ram_rdata<14> vdd 0.32fF
C8569 raven_soc_0|irq_pin BU_3VX2_47|Q 9.98fF
C8570 LS_3VX2_27|A vdd 3.91fF
C8571 raven_padframe_0|BT4F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C8572 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<11> 0.41fF
C8573 BU_3VX2_1|A vdd 0.18fF
C8574 BU_3VX2_12|A raven_soc_0|flash_io2_oeb 0.01fF
C8575 LS_3VX2_24|A LS_3VX2_16|A 0.01fF
C8576 raven_soc_0|gpio_pullup<0> BU_3VX2_24|Q 0.01fF
C8577 BU_3VX2_0|Q BU_3VX2_66|Q 0.01fF
C8578 raven_soc_0|gpio_outenb<1> BU_3VX2_26|Q 0.01fF
C8579 BU_3VX2_0|Q BU_3VX2_20|Q 0.01fF
C8580 VDD raven_padframe_0|VDDORPADF_3|GNDR 0.16fF
C8581 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<20> 33.18fF
C8582 raven_soc_0|ram_rdata<4> raven_soc_0|ram_addr<2> 0.31fF
C8583 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<10> 12.29fF
C8584 raven_soc_0|ram_rdata<30> raven_soc_0|ram_addr<3> 11.33fF
C8585 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<24> 2.18fF
C8586 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<31> 0.22fF
C8587 raven_soc_0|ram_rdata<8> raven_soc_0|ram_addr<4> 0.10fF
C8588 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_outenb<8> 3.23fF
C8589 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<6> 3.40fF
C8590 raven_soc_0|gpio_out<10> raven_soc_0|gpio_pullup<14> 0.01fF
C8591 BU_3VX2_37|Q BU_3VX2_32|Q 17.23fF
C8592 BU_3VX2_14|Q BU_3VX2_11|Q 13.54fF
C8593 raven_padframe_0|axtoc02_3v3_0|GNDR raven_padframe_0|axtoc02_3v3_0|GNDO 1.17fF
C8594 markings_0|manufacturer_0|_alphabet_L_0|m2_0_0# markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# 0.11fF
C8595 BU_3VX2_6|A BU_3VX2_12|A 1.89fF
C8596 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<11> 4.27fF
C8597 BU_3VX2_3|A raven_soc_0|flash_io2_do 0.01fF
C8598 BU_3VX2_23|A BU_3VX2_24|Q 0.03fF
C8599 LS_3VX2_3|Q raven_soc_0|flash_io2_di 0.01fF
C8600 BU_3VX2_15|A raven_soc_0|flash_io2_do 0.01fF
C8601 LS_3VX2_10|Q vdd 1.08fF
C8602 VDD raven_padframe_0|GNDORPADF_0|GNDOR 0.24fF
C8603 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<8> 1.10fF
C8604 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<10> 1.02fF
C8605 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<7> 0.15fF
C8606 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<11> 32.23fF
C8607 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<15> 0.43fF
C8608 BU_3VX2_0|Q raven_soc_0|ram_rdata<28> 0.02fF
C8609 BU_3VX2_24|A BU_3VX2_38|A 0.01fF
C8610 BU_3VX2_19|A BU_3VX2_28|A 2.34fF
C8611 BU_3VX2_18|A BU_3VX2_31|A 1.63fF
C8612 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<9> 0.01fF
C8613 LOGIC0_3V_4|Q raven_soc_0|flash_io2_di 0.08fF
C8614 BU_3VX2_65|A BU_3VX2_36|Q 0.03fF
C8615 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<13> 0.01fF
C8616 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<14> 215.78fF
C8617 raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<8> 0.59fF
C8618 raven_soc_0|gpio_out<1> BU_3VX2_40|Q 0.03fF
C8619 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<8> 1.23fF
C8620 raven_soc_0|gpio_out<12> raven_soc_0|gpio_outenb<9> 0.02fF
C8621 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pullup<14> 0.01fF
C8622 raven_soc_0|gpio_outenb<10> BU_3VX2_71|Q 0.01fF
C8623 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<14> 0.01fF
C8624 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<5> 0.01fF
C8625 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<1> 0.01fF
C8626 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<26> 0.06fF
C8627 BU_3VX2_6|Q BU_3VX2_38|Q 5.26fF
C8628 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<25> 25.10fF
C8629 BU_3VX2_19|Q BU_3VX2_2|Q 4.71fF
C8630 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<2> 6.13fF
C8631 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<19> 29.17fF
C8632 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<14> 0.17fF
C8633 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<13> 0.02fF
C8634 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<17> 6.74fF
C8635 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<21> 5.52fF
C8636 BU_3VX2_73|Q LS_3VX2_22|A 57.58fF
C8637 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<26> 9.93fF
C8638 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<22> 3.04fF
C8639 BU_3VX2_66|Q BU_3VX2_30|Q 6.73fF
C8640 BU_3VX2_2|Q BU_3VX2_18|Q 0.77fF
C8641 BU_3VX2_30|Q BU_3VX2_20|Q 7.34fF
C8642 BU_3VX2_19|Q BU_3VX2_10|Q 9.15fF
C8643 BU_3VX2_9|Q BU_3VX2_22|Q 4.24fF
C8644 BU_3VX2_18|Q BU_3VX2_10|Q 4.94fF
C8645 BU_3VX2_7|Q BU_3VX2_67|Q 0.07fF
C8646 BU_3VX2_6|Q BU_3VX2_67|Q 1.67fF
C8647 BU_3VX2_16|Q BU_3VX2_20|Q 9.17fF
C8648 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<13> 97.01fF
C8649 BU_3VX2_15|Q BU_3VX2_22|Q 4.66fF
C8650 BU_3VX2_69|Q BU_3VX2_17|Q 0.01fF
C8651 BU_3VX2_38|Q BU_3VX2_7|Q 4.36fF
C8652 raven_soc_0|gpio_pullup<5> vdd 1.06fF
C8653 BU_3VX2_54|A vdd 0.17fF
C8654 LS_3VX2_20|Q BU_3VX2_44|Q 0.63fF
C8655 LS_3VX2_12|A LS_3VX2_14|A 32.48fF
C8656 BU_3VX2_23|A BU_3VX2_13|A 2.11fF
C8657 raven_padframe_0|FILLER20F_7|VDDR raven_padframe_0|FILLER20F_7|GNDR 0.68fF
C8658 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<1> 9.34fF
C8659 raven_padframe_0|BBCUD4F_10|VDDO raven_padframe_0|BBCUD4F_10|GNDO 2.28fF
C8660 BU_3VX2_35|A BU_3VX2_0|Q 1.11fF
C8661 raven_padframe_0|aregc01_3v3_1|m4_0_31172# raven_padframe_0|aregc01_3v3_1|m4_0_30133# 0.02fF
C8662 BU_3VX2_17|A BU_3VX2_27|A 2.13fF
C8663 BU_3VX2_26|A raven_soc_0|flash_csb 5.53fF
C8664 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<11> 0.01fF
C8665 raven_soc_0|gpio_pulldown<15> BU_3VX2_0|Q 0.01fF
C8666 raven_padframe_0|axtoc02_3v3_0|m4_0_31172# raven_padframe_0|axtoc02_3v3_0|m4_0_30653# 0.17fF
C8667 BU_3VX2_63|Q raven_soc_0|gpio_pullup<3> 0.01fF
C8668 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<0> 0.01fF
C8669 LOGIC0_3V_1|Q LOGIC0_3V_0|Q 23.11fF
C8670 AMUX4_3V_3|SEL[1] BU_3VX2_23|Q 0.01fF
C8671 raven_soc_0|ram_addr<0> vdd 0.18fF
C8672 BU_3VX2_25|A BU_3VX2_5|A 0.01fF
C8673 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<15> 0.40fF
C8674 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<11> 0.01fF
C8675 BU_3VX2_11|A raven_soc_0|flash_csb 0.01fF
C8676 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<5> 0.07fF
C8677 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<2> 6.54fF
C8678 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<13> 1.76fF
C8679 raven_soc_0|gpio_out<7> raven_soc_0|gpio_out<11> 0.67fF
C8680 raven_padframe_0|BBCUD4F_1|VDDR raven_padframe_0|BBCUD4F_1|GNDR 0.68fF
C8681 markings_0|manufacturer_0|_alphabet_F_0|m2_0_0# markings_0|product_name_0|_alphabet_A_0|m2_0_0# 0.16fF
C8682 BU_3VX2_7|A raven_soc_0|flash_io3_do 0.01fF
C8683 VDD raven_padframe_0|FILLER20F_1|GNDO 0.07fF
C8684 raven_soc_0|gpio_outenb<3> raven_soc_0|ext_clk 0.01fF
C8685 BU_3VX2_31|A raven_soc_0|gpio_in<14> 0.01fF
C8686 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<5> 0.01fF
C8687 raven_soc_0|flash_io2_di raven_soc_0|flash_io1_oeb 20.05fF
C8688 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<15> 0.06fF
C8689 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<13> 0.20fF
C8690 BU_3VX2_1|Q AMUX4_3V_4|SEL[0] 0.93fF
C8691 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<16> 0.21fF
C8692 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<1> 1.68fF
C8693 raven_padframe_0|BBC4F_0|GNDR raven_padframe_0|BBC4F_0|VDDO 0.09fF
C8694 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<7> 0.37fF
C8695 raven_soc_0|gpio_in<1> BU_3VX2_26|Q 0.01fF
C8696 BU_3VX2_24|A BU_3VX2_23|Q 0.16fF
C8697 BU_3VX2_37|A BU_3VX2_35|Q 0.03fF
C8698 LS_3VX2_12|A BU_3VX2_56|Q 4.17fF
C8699 BU_3VX2_4|A raven_soc_0|flash_io0_di 0.07fF
C8700 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<12> 0.71fF
C8701 raven_padframe_0|BT4FC_0|VDDR raven_padframe_0|BT4FC_0|VDDO 0.06fF
C8702 LS_3VX2_8|A BU_3VX2_53|Q 6.77fF
C8703 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<13> 0.20fF
C8704 BU_3VX2_31|A raven_soc_0|gpio_pullup<6> 0.01fF
C8705 IN_3VX2_1|A BU_3VX2_24|Q 32.57fF
C8706 VDD raven_padframe_0|FILLER20F_2|VDDR 0.71fF
C8707 raven_soc_0|gpio_pullup<12> BU_3VX2_28|Q 0.01fF
C8708 raven_soc_0|gpio_outenb<12> vdd 0.27fF
C8709 VDD raven_padframe_0|FILLER20F_5|GNDO 0.07fF
C8710 LS_3VX2_13|A BU_3VX2_55|Q 0.01fF
C8711 raven_soc_0|gpio_pullup<11> apllc03_1v8_0|CLK 0.01fF
C8712 raven_soc_0|gpio_pullup<9> BU_3VX2_29|Q 0.01fF
C8713 BU_3VX2_38|A BU_3VX2_29|A 0.01fF
C8714 BU_3VX2_20|A BU_3VX2_26|A 3.62fF
C8715 BU_3VX2_12|A BU_3VX2_27|A 0.01fF
C8716 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<4> 0.02fF
C8717 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<12> 193.98fF
C8718 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<9> 1.90fF
C8719 LS_3VX2_3|A raven_soc_0|gpio_pullup<8> 0.01fF
C8720 BU_3VX2_35|A raven_soc_0|flash_io3_di 0.09fF
C8721 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<0> 0.01fF
C8722 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<22> 1.01fF
C8723 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<8> 14.26fF
C8724 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<7> 2.12fF
C8725 raven_soc_0|gpio_in<9> raven_soc_0|gpio_in<6> 1.94fF
C8726 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<11> 0.02fF
C8727 BU_3VX2_55|A LS_3VX2_17|Q 0.12fF
C8728 BU_3VX2_56|A LS_3VX2_16|Q 0.17fF
C8729 BU_3VX2_54|A BU_3VX2_62|A 0.15fF
C8730 BU_3VX2_57|A LS_3VX2_15|Q 0.27fF
C8731 BU_3VX2_58|A BU_3VX2_61|A 0.83fF
C8732 BU_3VX2_59|A BU_3VX2_60|A 5.87fF
C8733 raven_soc_0|gpio_in<10> VDD3V3 0.07fF
C8734 LS_3VX2_20|Q vdd 0.37fF
C8735 BU_3VX2_37|A BU_3VX2_38|A 33.57fF
C8736 BU_3VX2_32|A BU_3VX2_67|A 0.54fF
C8737 BU_3VX2_22|A BU_3VX2_18|A 5.07fF
C8738 raven_padframe_0|APR00DF_5|VDDR raven_padframe_0|APR00DF_5|GNDR 0.68fF
C8739 BU_3VX2_20|A BU_3VX2_11|A 1.75fF
C8740 BU_3VX2_71|A BU_3VX2_31|A 0.01fF
C8741 BU_3VX2_19|A BU_3VX2_14|A 3.76fF
C8742 raven_padframe_0|BBCUD4F_13|GNDR raven_padframe_0|BBCUD4F_13|VDDO 0.09fF
C8743 IN_3VX2_1|A BU_3VX2_13|A 0.01fF
C8744 raven_soc_0|gpio_pulldown<0> BU_3VX2_0|Q 0.01fF
C8745 BU_3VX2_31|A raven_soc_0|gpio_outenb<15> 0.01fF
C8746 raven_padframe_0|aregc01_3v3_0|m4_0_30653# raven_padframe_0|aregc01_3v3_0|m4_0_30133# 0.09fF
C8747 raven_padframe_0|aregc01_3v3_0|m4_0_31172# raven_padframe_0|aregc01_3v3_0|m4_0_29333# 0.01fF
C8748 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<12> 0.01fF
C8749 raven_padframe_0|BBCUD4F_0|GNDR raven_padframe_0|BBCUD4F_0|VDDO 0.09fF
C8750 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<4> 0.48fF
C8751 BU_3VX2_33|A raven_soc_0|gpio_pullup<15> 1.77fF
C8752 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<3> 1.37fF
C8753 markings_0|efabless_logo_0|m1_8700_n6150# markings_0|efabless_logo_0|m1_7500_n8250# 0.01fF
C8754 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<12> 73.89fF
C8755 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_pullup<5> 0.12fF
C8756 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<9> 22.79fF
C8757 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<14> 0.30fF
C8758 raven_soc_0|gpio_pullup<14> raven_soc_0|ext_clk 0.01fF
C8759 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<15> 0.02fF
C8760 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<13> 70.51fF
C8761 BU_3VX2_73|Q BU_3VX2_60|Q 0.01fF
C8762 BU_3VX2_10|Q BU_3VX2_27|Q 5.39fF
C8763 BU_3VX2_2|Q BU_3VX2_27|Q 19.17fF
C8764 BU_3VX2_1|Q vdd 1.71fF
C8765 raven_soc_0|ext_clk raven_padframe_0|ICF_2|PO 0.04fF
C8766 LS_3VX2_21|Q LS_3VX2_21|A 0.06fF
C8767 BU_3VX2_17|Q BU_3VX2_29|Q 2.87fF
C8768 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<2> 0.01fF
C8769 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<8> 0.01fF
C8770 IN_3VX2_1|Q VDD3V3 3.00fF
C8771 BU_3VX2_0|Q BU_3VX2_16|Q 0.01fF
C8772 VDD raven_padframe_0|APR00DF_3|GNDR 0.16fF
C8773 LS_3VX2_4|A BU_3VX2_53|Q 24.01fF
C8774 BU_3VX2_0|Q BU_3VX2_30|Q 0.12fF
C8775 VDD raven_padframe_0|FILLER02F_0|GNDR 0.20fF
C8776 raven_soc_0|ser_rx BU_3VX2_55|Q 1.68fF
C8777 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_out<8> 3.94fF
C8778 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<30> 0.25fF
C8779 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<24> 7.11fF
C8780 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<8> 10.74fF
C8781 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<4> 0.99fF
C8782 raven_soc_0|ram_rdata<22> raven_soc_0|ram_addr<4> 0.62fF
C8783 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<23> 0.01fF
C8784 raven_soc_0|flash_clk BU_3VX2_27|Q 10.25fF
C8785 raven_soc_0|ram_rdata<20> apllc03_1v8_0|CLK 0.01fF
C8786 markings_0|manufacturer_0|_alphabet_E_2|m2_0_0# markings_0|manufacturer_0|_alphabet_L_0|m2_0_0# 0.24fF
C8787 markings_0|product_name_0|_alphabet_1_0|m2_64_1376# markings_0|product_name_0|_alphabet_V_1|m2_0_560# 0.50fF
C8788 aopac01_3v3_0|IB VDD3V3 1.00fF
C8789 VDD raven_padframe_0|FILLER50F_1|GNDO 0.07fF
C8790 IN_3VX2_1|A raven_soc_0|gpio_out<15> 0.01fF
C8791 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<9> 0.69fF
C8792 raven_soc_0|gpio_in<0> VDD3V3 0.03fF
C8793 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<11> 23.16fF
C8794 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<9> 39.76fF
C8795 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<12> 0.03fF
C8796 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<13> 0.13fF
C8797 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<10> 0.09fF
C8798 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<14> 0.14fF
C8799 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<15> 0.34fF
C8800 raven_soc_0|gpio_out<11> BU_3VX2_40|Q 0.01fF
C8801 BU_3VX2_0|Q raven_soc_0|flash_io3_di 0.01fF
C8802 raven_soc_0|flash_csb VDD3V3 18.41fF
C8803 BU_3VX2_7|A BU_3VX2_8|A 24.20fF
C8804 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<13> 0.01fF
C8805 BU_3VX2_38|A LS_3VX2_3|Q 0.01fF
C8806 BU_3VX2_25|A BU_3VX2_24|Q 0.16fF
C8807 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<13> 0.99fF
C8808 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<8> 0.18fF
C8809 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<14> 14.07fF
C8810 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<8> 0.02fF
C8811 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<9> 1.19fF
C8812 raven_soc_0|gpio_pullup<10> BU_3VX2_71|Q 0.01fF
C8813 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pulldown<6> 0.02fF
C8814 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pullup<14> 0.01fF
C8815 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pullup<6> 3.78fF
C8816 raven_padframe_0|BBCUD4F_9|VDDR raven_padframe_0|BBCUD4F_9|VDDO 0.06fF
C8817 raven_soc_0|gpio_pulldown<8> apllc03_1v8_0|CLK 0.01fF
C8818 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<28> 7.86fF
C8819 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<27> 0.64fF
C8820 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<29> 0.67fF
C8821 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<26> 0.08fF
C8822 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<3> 0.02fF
C8823 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<1> 0.11fF
C8824 BU_3VX2_13|Q BU_3VX2_68|Q 35.03fF
C8825 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<13> 31.03fF
C8826 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<14> 33.30fF
C8827 BU_3VX2_12|Q BU_3VX2_5|Q 5.10fF
C8828 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<2> 1.64fF
C8829 BU_3VX2_35|Q BU_3VX2_38|Q 53.84fF
C8830 BU_3VX2_65|Q BU_3VX2_7|Q 0.08fF
C8831 BU_3VX2_64|Q BU_3VX2_22|Q 1.03fF
C8832 BU_3VX2_43|A BU_3VX2_43|Q 0.10fF
C8833 AMUX4_3V_0|SEL[0] LS_3VX2_20|A 7.50fF
C8834 raven_padframe_0|CORNERESDF_3|VDDR raven_padframe_0|CORNERESDF_3|GNDO 0.13fF
C8835 LS_3VX2_9|A LS_3VX2_11|A 23.36fF
C8836 BU_3VX2_35|A BU_3VX2_63|A 0.08fF
C8837 BU_3VX2_21|A BU_3VX2_18|A 7.13fF
C8838 BU_3VX2_5|A BU_3VX2_4|A 21.57fF
C8839 LS_3VX2_9|Q LS_3VX2_5|A 0.54fF
C8840 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<11> 13.01fF
C8841 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<10> 1.07fF
C8842 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<5> 0.01fF
C8843 raven_soc_0|ram_addr<9> vdd 0.16fF
C8844 raven_soc_0|ram_wdata<29> vdd 1.96fF
C8845 BU_3VX2_56|Q BU_3VX2_46|Q 0.10fF
C8846 raven_soc_0|ram_wdata<17> apllc03_1v8_0|CLK 0.01fF
C8847 BU_3VX2_22|A BU_3VX2_71|A 0.02fF
C8848 LS_3VX2_11|Q LS_3VX2_8|A 0.18fF
C8849 BU_3VX2_25|A BU_3VX2_13|A 1.75fF
C8850 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<14> 0.47fF
C8851 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<6> 0.01fF
C8852 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<11> 0.01fF
C8853 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<13> 9.61fF
C8854 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<12> 8.82fF
C8855 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<6> 0.01fF
C8856 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<11> 0.02fF
C8857 markings_0|efabless_logo_0|m1_3300_n1350# markings_0|efabless_logo_0|m1_2400_n2250# 0.25fF
C8858 BU_3VX2_38|A BU_3VX2_38|Q 0.08fF
C8859 BU_3VX2_20|A VDD3V3 0.43fF
C8860 BU_3VX2_1|Q BU_3VX2_70|Q 0.55fF
C8861 raven_soc_0|ram_rdata<24> raven_soc_0|ram_addr<0> 6.91fF
C8862 raven_soc_0|flash_io1_di raven_soc_0|flash_io0_do 40.98fF
C8863 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<15> 19.86fF
C8864 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<13> 7.57fF
C8865 raven_soc_0|flash_io0_oeb raven_soc_0|flash_io0_di 16.95fF
C8866 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<29> 3.31fF
C8867 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<27> 0.01fF
C8868 raven_soc_0|flash_io2_oeb raven_soc_0|flash_clk 78.16fF
C8869 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<31> 7.52fF
C8870 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<17> 0.01fF
C8871 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<24> 0.01fF
C8872 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<16> 2.20fF
C8873 markings_0|date_0|_alphabet_8_0|m2_9_235# markings_0|date_0|_alphabet_1_1|m2_64_1376# 0.36fF
C8874 raven_padframe_0|FILLER20F_2|VDDR raven_padframe_0|FILLER20F_2|GNDO 0.13fF
C8875 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<9> 0.01fF
C8876 BU_3VX2_6|A raven_soc_0|flash_clk 0.01fF
C8877 LS_3VX2_22|Q LS_3VX2_22|A 0.05fF
C8878 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<5> 0.54fF
C8879 BU_3VX2_38|A raven_soc_0|flash_io1_oeb 0.01fF
C8880 BU_3VX2_9|A raven_soc_0|flash_io2_oeb 0.01fF
C8881 BU_3VX2_19|A raven_soc_0|flash_io1_do 0.01fF
C8882 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<13> 5.44fF
C8883 LS_3VX2_7|A adc0_data<5> 0.06fF
C8884 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<6> 0.08fF
C8885 VDD raven_padframe_0|aregc01_3v3_0|GNDO 0.06fF
C8886 VDD raven_padframe_0|CORNERESDF_0|GNDR 0.16fF
C8887 BU_3VX2_28|A BU_3VX2_27|Q 0.16fF
C8888 LS_3VX2_13|A BU_3VX2_57|Q 0.01fF
C8889 raven_soc_0|gpio_outenb<0> BU_3VX2_28|Q 0.01fF
C8890 raven_soc_0|gpio_pulldown<9> BU_3VX2_29|Q 0.01fF
C8891 VDD raven_padframe_0|BBCUD4F_2|GNDO 0.07fF
C8892 raven_soc_0|gpio_pullup<12> vdd 0.24fF
C8893 BU_3VX2_6|A BU_3VX2_9|A 4.74fF
C8894 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<0> 0.01fF
C8895 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<7> 0.01fF
C8896 BU_3VX2_63|Q raven_soc_0|flash_io0_oeb 0.01fF
C8897 BU_3VX2_40|Q raven_soc_0|gpio_in<12> 0.01fF
C8898 raven_soc_0|ext_clk raven_soc_0|gpio_in<9> 0.01fF
C8899 BU_3VX2_52|A BU_3VX2_57|A 0.96fF
C8900 BU_3VX2_54|A BU_3VX2_55|A 11.16fF
C8901 BU_3VX2_53|A BU_3VX2_56|A 1.94fF
C8902 VDD3V3 BU_3VX2_59|A 0.05fF
C8903 BU_3VX2_24|A BU_3VX2_31|A 5.26fF
C8904 raven_soc_0|gpio_in<13> VDD3V3 0.07fF
C8905 raven_spi_0|SDO raven_soc_0|gpio_pulldown<15> 1.30fF
C8906 BU_3VX2_1|A BU_3VX2_69|A 0.54fF
C8907 LOGIC0_3V_4|Q raven_soc_0|gpio_out<4> 0.01fF
C8908 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_in<3> 1.22fF
C8909 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<10> 0.02fF
C8910 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<5> 0.01fF
C8911 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<12> 0.01fF
C8912 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<14> 0.06fF
C8913 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<8> 28.02fF
C8914 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<23> 0.02fF
C8915 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<19> 0.27fF
C8916 raven_soc_0|flash_io3_di raven_soc_0|irq_pin 0.01fF
C8917 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<14> 0.02fF
C8918 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<7> 49.85fF
C8919 BU_3VX2_38|Q BU_3VX2_23|Q 0.26fF
C8920 BU_3VX2_12|Q BU_3VX2_28|Q 1.86fF
C8921 BU_3VX2_13|Q BU_3VX2_24|Q 4.65fF
C8922 BU_3VX2_2|Q BU_3VX2_25|Q 7.19fF
C8923 BU_3VX2_66|Q BU_3VX2_26|Q 0.97fF
C8924 BU_3VX2_73|Q BU_3VX2_62|Q 0.01fF
C8925 BU_3VX2_15|Q apllc03_1v8_0|CLK 0.01fF
C8926 BU_3VX2_10|Q BU_3VX2_25|Q 2.60fF
C8927 BU_3VX2_67|Q BU_3VX2_23|Q 2.81fF
C8928 BU_3VX2_20|Q BU_3VX2_26|Q 6.06fF
C8929 LS_3VX2_21|Q LS_3VX2_27|A 0.20fF
C8930 BU_3VX2_9|Q apllc03_1v8_0|CLK 0.01fF
C8931 BU_3VX2_53|Q vdd 1.87fF
C8932 BU_3VX2_55|Q BU_3VX2_72|Q 1.07fF
C8933 raven_spi_0|CSB BU_3VX2_33|A 35.89fF
C8934 BU_3VX2_21|A BU_3VX2_71|A 0.01fF
C8935 raven_padframe_0|VDDPADFC_0|VDDR LOGIC0_3V_4|Q 0.01fF
C8936 BU_3VX2_32|A BU_3VX2_33|Q 0.03fF
C8937 LS_3VX2_5|A BU_3VX2_73|Q 7.26fF
C8938 raven_soc_0|ser_rx BU_3VX2_57|Q 2.01fF
C8939 BU_3VX2_0|Q AMUX4_3V_3|SEL[0] 12.66fF
C8940 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pullup<6> 51.33fF
C8941 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<10> 1.15fF
C8942 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<5> 3.11fF
C8943 raven_soc_0|ram_rdata<13> raven_soc_0|ram_rdata<16> 17.95fF
C8944 BU_3VX2_47|A vdd 0.06fF
C8945 raven_soc_0|flash_clk BU_3VX2_25|Q 0.01fF
C8946 raven_soc_0|flash_io0_di BU_3VX2_29|Q 0.01fF
C8947 AMUX4_3V_0|SEL[0] BU_3VX2_47|Q 13.03fF
C8948 raven_soc_0|flash_io1_oeb BU_3VX2_23|Q 0.01fF
C8949 raven_soc_0|flash_io0_do BU_3VX2_28|Q 0.01fF
C8950 raven_padframe_0|FILLER50F_0|GNDR raven_padframe_0|FILLER50F_0|GNDO 0.81fF
C8951 raven_padframe_0|aregc01_3v3_1|GNDR raven_padframe_0|aregc01_3v3_1|GNDO 0.59fF
C8952 markings_0|manufacturer_0|_alphabet_S_1|m2_32_224# markings_0|manufacturer_0|_alphabet_E_2|m2_0_0# 0.01fF
C8953 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<8> 0.14fF
C8954 BU_3VX2_10|A raven_soc_0|flash_io0_do 0.03fF
C8955 LS_3VX2_10|A LS_3VX2_19|A 0.01fF
C8956 LS_3VX2_10|A BU_3VX2_52|Q 15.01fF
C8957 BU_3VX2_63|A raven_soc_0|flash_io3_di 0.01fF
C8958 BU_3VX2_13|A BU_3VX2_13|Q 0.08fF
C8959 BU_3VX2_28|A raven_soc_0|flash_io2_oeb 5.83fF
C8960 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<14> 0.56fF
C8961 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<9> 15.76fF
C8962 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<12> 0.02fF
C8963 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<10> 6.11fF
C8964 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<15> 0.02fF
C8965 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<11> 12.57fF
C8966 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<13> 0.02fF
C8967 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pullup<5> 0.02fF
C8968 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<11> 0.02fF
C8969 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<20> 1.12fF
C8970 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<0> 1.32fF
C8971 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<23> 3.98fF
C8972 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<19> 0.02fF
C8973 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<28> 0.02fF
C8974 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<13> 0.01fF
C8975 BU_3VX2_6|A BU_3VX2_28|A 0.01fF
C8976 BU_3VX2_5|A raven_soc_0|flash_io0_oeb 0.01fF
C8977 BU_3VX2_0|A raven_soc_0|flash_io0_do 5.07fF
C8978 IN_3VX2_1|A raven_soc_0|gpio_out<10> 0.01fF
C8979 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_pullup<13> 0.04fF
C8980 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<9> 0.02fF
C8981 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pullup<14> 1.04fF
C8982 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<29> 0.04fF
C8983 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<13> 0.05fF
C8984 raven_soc_0|gpio_pulldown<4> BU_3VX2_71|Q 0.01fF
C8985 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pulldown<7> 10.45fF
C8986 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pulldown<6> 0.02fF
C8987 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pullup<6> 0.02fF
C8988 BU_3VX2_27|A raven_soc_0|flash_clk 8.01fF
C8989 LS_3VX2_13|A LS_3VX2_16|A 0.01fF
C8990 raven_soc_0|gpio_pulldown<15> BU_3VX2_26|Q 0.01fF
C8991 raven_soc_0|gpio_pulldown<14> BU_3VX2_28|Q 0.01fF
C8992 BU_3VX2_63|Q BU_3VX2_29|Q 2.83fF
C8993 raven_padframe_0|BBCUD4F_2|VDDR raven_padframe_0|BBCUD4F_2|GNDO 0.13fF
C8994 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<12> 86.85fF
C8995 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<12> 0.02fF
C8996 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<2> 13.96fF
C8997 BU_3VX2_68|Q BU_3VX2_69|Q 27.68fF
C8998 BU_3VX2_64|Q BU_3VX2_31|Q 1.26fF
C8999 AMUX4_3V_4|SEL[1] BU_3VX2_33|Q 9.42fF
C9000 BU_3VX2_44|A BU_3VX2_42|Q 0.03fF
C9001 raven_padframe_0|FILLER40F_0|GNDR raven_padframe_0|FILLER40F_0|GNDO 0.81fF
C9002 raven_padframe_0|CORNERESDF_2|GNDR raven_padframe_0|CORNERESDF_2|GNDO 0.81fF
C9003 BU_3VX2_9|A BU_3VX2_27|A 0.01fF
C9004 BU_3VX2_16|A BU_3VX2_31|A 0.01fF
C9005 BU_3VX2_4|A BU_3VX2_13|A 1.14fF
C9006 BU_3VX2_31|A BU_3VX2_29|A 31.12fF
C9007 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pulldown<12> 14.26fF
C9008 BU_3VX2_24|A BU_3VX2_22|A 13.39fF
C9009 raven_soc_0|flash_io2_oeb BU_3VX2_33|Q 0.01fF
C9010 raven_soc_0|ram_rdata<29> vdd 0.27fF
C9011 BU_3VX2_73|Q BU_3VX2_45|Q 7.18fF
C9012 raven_soc_0|ram_wdata<18> apllc03_1v8_0|CLK 0.01fF
C9013 AMUX4_3V_1|SEL[0] BU_3VX2_55|Q 26.38fF
C9014 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<5> 0.01fF
C9015 BU_3VX2_37|A BU_3VX2_31|A 0.01fF
C9016 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<15> 0.01fF
C9017 BU_3VX2_67|A BU_3VX2_64|A 4.79fF
C9018 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_out<3> 2.95fF
C9019 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<2> 1.69fF
C9020 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<8> 0.01fF
C9021 IN_3VX2_1|A raven_soc_0|gpio_out<9> 0.01fF
C9022 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<5> 1.97fF
C9023 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_outenb<15> 1.08fF
C9024 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<14> 12.67fF
C9025 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<12> 0.01fF
C9026 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<13> 15.86fF
C9027 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<11> 11.09fF
C9028 raven_soc_0|gpio_pullup<0> raven_soc_0|ext_clk 0.01fF
C9029 raven_soc_0|gpio_outenb<1> VDD3V3 1.65fF
C9030 adc_high BU_3VX2_52|A 0.02fF
C9031 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<6> 1.05fF
C9032 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<31> 19.61fF
C9033 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<9> 1.22fF
C9034 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<3> 18.29fF
C9035 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<6> 0.01fF
C9036 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<24> 0.01fF
C9037 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<23> 0.01fF
C9038 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<20> 0.01fF
C9039 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<13> 5.35fF
C9040 BU_3VX2_6|Q BU_3VX2_36|Q 13.82fF
C9041 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<26> 0.02fF
C9042 raven_soc_0|flash_io2_do raven_soc_0|flash_io0_di 45.77fF
C9043 BU_3VX2_4|Q BU_3VX2_67|Q 1.31fF
C9044 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<1> 0.15fF
C9045 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<2> 2.17fF
C9046 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<27> 0.02fF
C9047 BU_3VX2_36|Q BU_3VX2_7|Q 0.44fF
C9048 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<19> 144.39fF
C9049 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<22> 159.15fF
C9050 BU_3VX2_38|Q BU_3VX2_4|Q 8.90fF
C9051 raven_soc_0|ram_rdata<31> raven_soc_0|ram_wdata<13> 0.01fF
C9052 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<29> 0.01fF
C9053 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<17> 3.52fF
C9054 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<31> 0.01fF
C9055 BU_3VX2_11|Q BU_3VX2_20|Q 3.52fF
C9056 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<21> 0.01fF
C9057 AMUX4_3V_0|SEL[1] BU_3VX2_59|Q 1.34fF
C9058 LOGIC0_3V_0|Q LOGIC0_3V_2|Q 7.53fF
C9059 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<9> 0.01fF
C9060 raven_spi_0|SDO raven_soc_0|flash_io3_di 0.84fF
C9061 BU_3VX2_23|A raven_soc_0|ext_clk 0.01fF
C9062 VDD raven_padframe_0|ICF_1|GNDR 0.16fF
C9063 BU_3VX2_28|A BU_3VX2_25|Q 0.02fF
C9064 raven_soc_0|gpio_pulldown<13> BU_3VX2_23|Q 0.01fF
C9065 raven_soc_0|ser_rx LS_3VX2_16|A 7.06fF
C9066 raven_soc_0|gpio_pulldown<10> BU_3VX2_28|Q 0.01fF
C9067 raven_soc_0|gpio_outenb<0> vdd 0.20fF
C9068 BU_3VX2_0|Q BU_3VX2_26|Q 0.02fF
C9069 LS_3VX2_3|A BU_3VX2_27|Q 0.01fF
C9070 BU_3VX2_71|Q raven_soc_0|flash_io2_di 0.02fF
C9071 LS_3VX2_6|Q LS_3VX2_7|A 0.16fF
C9072 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<13> 0.01fF
C9073 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pulldown<10> 10.96fF
C9074 LS_3VX2_10|A BU_3VX2_58|Q 7.43fF
C9075 IN_3VX2_1|Q adc0_data<5> 0.77fF
C9076 VDD raven_padframe_0|BBC4F_2|GNDR 0.16fF
C9077 LS_3VX2_11|Q vdd 0.99fF
C9078 BU_3VX2_14|A raven_soc_0|flash_io2_oeb 0.01fF
C9079 BU_3VX2_63|Q raven_soc_0|flash_io2_do 0.01fF
C9080 raven_soc_0|gpio_pulldown<0> BU_3VX2_26|Q 0.01fF
C9081 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<15> 0.02fF
C9082 raven_soc_0|gpio_pullup<1> BU_3VX2_23|Q 0.01fF
C9083 raven_soc_0|gpio_outenb<2> apllc03_1v8_0|CLK 0.01fF
C9084 raven_soc_0|gpio_out<2> BU_3VX2_29|Q 0.01fF
C9085 AMUX4_3V_1|AOUT VDD3V3 8.49fF
C9086 BU_3VX2_43|A LS_3VX2_27|Q 0.82fF
C9087 BU_3VX2_44|A BU_3VX2_42|A 0.73fF
C9088 LS_3VX2_20|Q LS_3VX2_21|Q 16.46fF
C9089 VDD3V3 LS_3VX2_20|A 0.43fF
C9090 BU_3VX2_6|A BU_3VX2_14|A 1.39fF
C9091 LS_3VX2_3|Q BU_3VX2_31|A 0.01fF
C9092 BU_3VX2_28|A BU_3VX2_27|A 86.18fF
C9093 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<6> 0.63fF
C9094 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<4> 11.10fF
C9095 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<1> 0.61fF
C9096 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<0> 5.34fF
C9097 markings_0|efabless_logo_0|m1_2400_n2250# markings_0|efabless_logo_0|m1_1500_n3150# 0.19fF
C9098 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<13> 9.53fF
C9099 raven_soc_0|gpio_pulldown<11> BU_3VX2_71|Q 0.01fF
C9100 BU_3VX2_24|A BU_3VX2_21|A 7.80fF
C9101 raven_soc_0|gpio_pulldown<7> BU_3VX2_40|Q 0.30fF
C9102 raven_soc_0|gpio_pulldown<3> VDD3V3 0.22fF
C9103 BU_3VX2_12|Q vdd 0.83fF
C9104 LS_3VX2_22|A BU_3VX2_50|Q 6.95fF
C9105 BU_3VX2_16|Q BU_3VX2_26|Q 3.51fF
C9106 BU_3VX2_30|Q BU_3VX2_26|Q 9.71fF
C9107 BU_3VX2_69|Q BU_3VX2_24|Q 1.56fF
C9108 BU_3VX2_5|Q BU_3VX2_28|Q 0.31fF
C9109 LS_3VX2_17|A BU_3VX2_55|Q 9.52fF
C9110 BU_3VX2_68|Q BU_3VX2_29|Q 0.85fF
C9111 BU_3VX2_65|Q BU_3VX2_23|Q 0.32fF
C9112 BU_3VX2_57|Q BU_3VX2_72|Q 0.16fF
C9113 BU_3VX2_64|Q apllc03_1v8_0|CLK 0.98fF
C9114 BU_3VX2_22|A BU_3VX2_16|A 3.03fF
C9115 VDD raven_padframe_0|FILLER02F_0|VDDR 0.71fF
C9116 BU_3VX2_3|A BU_3VX2_17|A 0.01fF
C9117 BU_3VX2_22|A BU_3VX2_29|A 3.09fF
C9118 LOGIC1_3V_1|Q LOGIC0_3V_3|Q 0.32fF
C9119 BU_3VX2_15|A BU_3VX2_17|A 14.01fF
C9120 BU_3VX2_67|A BU_3VX2_66|A 24.87fF
C9121 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<12> 0.09fF
C9122 BU_3VX2_19|A raven_soc_0|flash_csb 1.59fF
C9123 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<4> 1.16fF
C9124 BU_3VX2_1|Q LS_3VX2_2|A 2.83fF
C9125 LS_3VX2_19|A raven_soc_0|ser_tx 103.66fF
C9126 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<16> 0.01fF
C9127 raven_soc_0|ram_wdata<31> raven_soc_0|ram_rdata<17> 1.04fF
C9128 raven_soc_0|ram_wdata<27> raven_soc_0|ram_addr<0> 0.01fF
C9129 raven_soc_0|flash_io0_do vdd 6.24fF
C9130 raven_soc_0|flash_io0_oeb BU_3VX2_24|Q 0.01fF
C9131 raven_soc_0|flash_io3_di BU_3VX2_26|Q 0.01fF
C9132 raven_soc_0|flash_io1_do BU_3VX2_27|Q 0.01fF
C9133 raven_soc_0|flash_io1_di BU_3VX2_28|Q 0.01fF
C9134 BU_3VX2_56|A BU_3VX2_58|Q 0.04fF
C9135 raven_padframe_0|FILLER01F_1|VDDR raven_padframe_0|FILLER01F_1|GNDR 0.68fF
C9136 raven_padframe_0|BT4FC_0|VDDO raven_padframe_0|BT4FC_0|GNDO 2.28fF
C9137 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<3> 1.04fF
C9138 raven_padframe_0|FILLER01F_0|GNDR raven_padframe_0|FILLER01F_0|GNDO 0.81fF
C9139 raven_padframe_0|FILLER02F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C9140 raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# raven_padframe_0|axtoc02_3v3_0|m4_55000_22024# 0.03fF
C9141 raven_padframe_0|axtoc02_3v3_0|m4_0_29333# raven_padframe_0|axtoc02_3v3_0|GNDO 0.25fF
C9142 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<13> 0.02fF
C9143 raven_soc_0|gpio_in<1> VDD3V3 1.85fF
C9144 BU_3VX2_10|A raven_soc_0|flash_io1_di 0.05fF
C9145 LS_3VX2_19|Q LS_3VX2_19|A 0.05fF
C9146 LS_3VX2_10|A LS_3VX2_22|A 11.15fF
C9147 BU_3VX2_20|A BU_3VX2_21|Q 0.03fF
C9148 IN_3VX2_1|A raven_soc_0|ext_clk 0.12fF
C9149 LS_3VX2_24|A LS_3VX2_19|A 1.23fF
C9150 LS_3VX2_24|A BU_3VX2_52|Q 0.02fF
C9151 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<12> 4.80fF
C9152 LS_3VX2_3|A raven_soc_0|flash_io2_oeb 0.05fF
C9153 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<8> 12.63fF
C9154 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<9> 8.40fF
C9155 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<15> 0.02fF
C9156 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<13> 0.02fF
C9157 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pullup<5> 0.02fF
C9158 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<14> 6.97fF
C9159 raven_soc_0|gpio_outenb<5> VDD3V3 0.11fF
C9160 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<0> 1.53fF
C9161 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<28> 7.67fF
C9162 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<19> 128.32fF
C9163 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<20> 0.12fF
C9164 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<23> 0.12fF
C9165 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<11> 13.38fF
C9166 raven_soc_0|gpio_out<1> BU_3VX2_63|Q 0.01fF
C9167 BU_3VX2_0|A raven_soc_0|flash_io1_di 17.03fF
C9168 BU_3VX2_40|A raven_soc_0|flash_io0_do 0.01fF
C9169 BU_3VX2_5|A raven_soc_0|flash_io2_do 0.01fF
C9170 BU_3VX2_31|A raven_soc_0|flash_io1_oeb 30.83fF
C9171 BU_3VX2_13|A raven_soc_0|flash_io0_oeb 0.01fF
C9172 adc_low raven_soc_0|ser_tx 0.05fF
C9173 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<5> 0.81fF
C9174 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<6> 0.82fF
C9175 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<9> 0.01fF
C9176 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<3> 0.02fF
C9177 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<14> 0.43fF
C9178 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<13> 0.59fF
C9179 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pulldown<7> 19.48fF
C9180 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<14> 0.01fF
C9181 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<15> 2.04fF
C9182 BU_3VX2_0|Q BU_3VX2_11|Q 0.01fF
C9183 BU_3VX2_33|A raven_soc_0|flash_io3_oeb 0.18fF
C9184 BU_3VX2_0|Q raven_soc_0|gpio_outenb<13> 0.01fF
C9185 VDD raven_padframe_0|axtoc02_3v3_0|GNDR 0.20fF
C9186 raven_soc_0|gpio_pulldown<14> vdd 0.15fF
C9187 AMUX2_3V_0|SEL BU_3VX2_51|Q 6.92fF
C9188 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<0> 4.97fF
C9189 BU_3VX2_20|A BU_3VX2_19|A 37.24fF
C9190 BU_3VX2_3|A BU_3VX2_12|A 1.10fF
C9191 BU_3VX2_68|A BU_3VX2_65|A 4.82fF
C9192 BU_3VX2_15|A BU_3VX2_12|A 7.02fF
C9193 LS_3VX2_8|A LS_3VX2_4|A 10.79fF
C9194 LS_3VX2_24|A adc_low 0.13fF
C9195 LOGIC0_3V_4|Q raven_soc_0|gpio_out<8> 0.01fF
C9196 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<8> 0.38fF
C9197 raven_padframe_0|BT4F_0|VDDR raven_padframe_0|BT4F_0|GNDR 0.68fF
C9198 BU_3VX2_73|Q AMUX4_3V_4|AIN3 0.02fF
C9199 raven_soc_0|ram_rdata<25> vdd 0.81fF
C9200 AMUX4_3V_1|SEL[0] BU_3VX2_57|Q 16.83fF
C9201 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<6> 0.01fF
C9202 BU_3VX2_22|A LS_3VX2_3|Q 0.77fF
C9203 BU_3VX2_21|A BU_3VX2_16|A 3.74fF
C9204 BU_3VX2_21|A BU_3VX2_29|A 2.63fF
C9205 BU_3VX2_14|A BU_3VX2_27|A 1.54fF
C9206 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<14> 0.01fF
C9207 IN_3VX2_1|A raven_soc_0|gpio_outenb<10> 0.01fF
C9208 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<11> 0.01fF
C9209 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<12> 0.01fF
C9210 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<6> 4.25fF
C9211 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<14> 15.97fF
C9212 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_outenb<15> 0.03fF
C9213 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<3> 7.50fF
C9214 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<11> 9.32fF
C9215 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<5> 0.01fF
C9216 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<9> 3.28fF
C9217 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<31> 0.01fF
C9218 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<24> 18.95fF
C9219 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<30> 25.89fF
C9220 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<23> 0.05fF
C9221 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<14> 0.18fF
C9222 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<21> 0.09fF
C9223 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<24> 9.31fF
C9224 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<20> 8.33fF
C9225 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<22> 0.01fF
C9226 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<7> 3.17fF
C9227 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<2> 3.74fF
C9228 raven_soc_0|flash_io1_do raven_soc_0|flash_io2_oeb 91.69fF
C9229 BU_3VX2_16|Q BU_3VX2_11|Q 15.80fF
C9230 BU_3VX2_14|Q BU_3VX2_8|Q 6.41fF
C9231 BU_3VX2_3|Q BU_3VX2_67|Q 2.90fF
C9232 BU_3VX2_21|Q BU_3VX2_14|Q 11.26fF
C9233 BU_3VX2_4|Q BU_3VX2_65|Q 6.79fF
C9234 raven_soc_0|flash_io3_do raven_soc_0|flash_io3_oeb 54.46fF
C9235 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<17> 0.02fF
C9236 BU_3VX2_12|Q BU_3VX2_70|Q 0.13fF
C9237 BU_3VX2_38|Q BU_3VX2_3|Q 12.33fF
C9238 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<21> 2.91fF
C9239 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<26> 0.06fF
C9240 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<8> 68.99fF
C9241 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<25> 0.15fF
C9242 BU_3VX2_2|Q BU_3VX2_37|Q 71.24fF
C9243 BU_3VX2_37|Q BU_3VX2_10|Q 3.89fF
C9244 VDD3V3 BU_3VX2_47|Q 0.02fF
C9245 BU_3VX2_24|Q BU_3VX2_29|Q 52.56fF
C9246 BU_3VX2_25|Q apllc03_1v8_0|B_CP 0.97fF
C9247 apllc03_1v8_0|B_VCO apllc03_1v8_0|CLK 3.93fF
C9248 LOGIC0_3V_4|Q raven_soc_0|gpio_out<6> 0.01fF
C9249 BU_3VX2_6|A raven_soc_0|flash_io1_do 0.02fF
C9250 BU_3VX2_2|A raven_soc_0|flash_io3_do 0.02fF
C9251 LOGIC1_3V_1|Q VDD3V3 0.06fF
C9252 LS_3VX2_11|A BU_3VX2_73|Q 9.62fF
C9253 BU_3VX2_64|A BU_3VX2_33|Q 0.02fF
C9254 LS_3VX2_3|A BU_3VX2_25|Q 0.01fF
C9255 VDD raven_padframe_0|aregc01_3v3_0|m4_0_31172# 0.12fF
C9256 raven_soc_0|gpio_pulldown<10> vdd 0.14fF
C9257 raven_soc_0|gpio_pulldown<12> BU_3VX2_28|Q 0.01fF
C9258 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<15> 11.05fF
C9259 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<13> 7.02fF
C9260 raven_soc_0|ram_rdata<0> raven_soc_0|ram_addr<0> 1.29fF
C9261 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<16> 10.15fF
C9262 raven_soc_0|ser_tx BU_3VX2_58|Q 7.50fF
C9263 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<2> 18.91fF
C9264 BU_3VX2_25|A raven_soc_0|ext_clk 0.01fF
C9265 LS_3VX2_10|A BU_3VX2_60|Q 0.01fF
C9266 LS_3VX2_24|A BU_3VX2_58|Q 0.01fF
C9267 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<5> 0.01fF
C9268 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<14> 0.02fF
C9269 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<8> 0.01fF
C9270 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<11> 0.01fF
C9271 BU_3VX2_10|A BU_3VX2_0|A 0.15fF
C9272 BU_3VX2_31|A raven_soc_0|gpio_pulldown<13> 0.01fF
C9273 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<10> 0.08fF
C9274 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<8> 7.55fF
C9275 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<10> 0.01fF
C9276 BU_3VX2_70|A BU_3VX2_33|A 0.96fF
C9277 BU_3VX2_22|A raven_soc_0|flash_io1_oeb 1.62fF
C9278 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<14> 0.03fF
C9279 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<6> 3.32fF
C9280 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<13> 14.18fF
C9281 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<14> 0.02fF
C9282 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<9> 0.01fF
C9283 raven_soc_0|gpio_out<11> raven_soc_0|flash_io0_di 0.01fF
C9284 BU_3VX2_5|Q vdd 1.19fF
C9285 LS_3VX2_17|A BU_3VX2_57|Q 12.05fF
C9286 LS_3VX2_22|A BU_3VX2_48|Q 5.65fF
C9287 VDD3V3 raven_padframe_0|VDDPADFC_0|GNDO 0.07fF
C9288 BU_3VX2_21|A LS_3VX2_3|Q 0.02fF
C9289 LS_3VX2_13|Q LS_3VX2_13|A 0.05fF
C9290 BU_3VX2_35|A BU_3VX2_26|A 0.28fF
C9291 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<0> 4.02fF
C9292 BU_3VX2_31|A raven_soc_0|gpio_pullup<1> 0.01fF
C9293 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<2> 0.10fF
C9294 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<0> 93.67fF
C9295 LS_3VX2_22|A raven_soc_0|ser_tx 0.01fF
C9296 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<27> 0.01fF
C9297 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<31> 0.01fF
C9298 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<17> 0.01fF
C9299 raven_soc_0|ram_wdata<17> raven_soc_0|ram_rdata<15> 0.01fF
C9300 raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<16> 0.06fF
C9301 raven_soc_0|ram_wdata<29> raven_soc_0|ram_wdata<27> 73.05fF
C9302 BU_3VX2_73|Q LS_3VX2_21|A 34.49fF
C9303 raven_soc_0|ram_wdata<22> raven_soc_0|ram_wdata<31> 10.27fF
C9304 raven_soc_0|ram_wdata<26> raven_soc_0|ram_addr<0> 0.01fF
C9305 raven_soc_0|ram_wdata<21> raven_soc_0|ram_rdata<13> 0.01fF
C9306 raven_soc_0|ram_wdata<25> raven_soc_0|ram_rdata<1> 2.09fF
C9307 raven_soc_0|ram_wdata<19> raven_soc_0|ram_rdata<17> 0.01fF
C9308 raven_soc_0|gpio_in<10> BU_3VX2_27|Q 0.01fF
C9309 raven_soc_0|flash_io1_di vdd 2.56fF
C9310 BU_3VX2_48|A BU_3VX2_42|A 0.16fF
C9311 BU_3VX2_47|A LS_3VX2_21|Q 0.17fF
C9312 BU_3VX2_41|A BU_3VX2_43|A 0.60fF
C9313 BU_3VX2_61|A BU_3VX2_61|Q 0.10fF
C9314 raven_soc_0|flash_io2_do BU_3VX2_24|Q 0.01fF
C9315 AMUX4_3V_1|SEL[0] LS_3VX2_16|A 7.54fF
C9316 raven_soc_0|flash_io3_do apllc03_1v8_0|CLK 13.78fF
C9317 raven_soc_0|flash_io1_do BU_3VX2_25|Q 0.01fF
C9318 raven_soc_0|gpio_out<15> BU_3VX2_29|Q 0.01fF
C9319 BU_3VX2_35|A BU_3VX2_11|A 1.74fF
C9320 BU_3VX2_35|A LOGIC0_3V_3|Q 0.04fF
C9321 raven_padframe_0|aregc01_3v3_1|m4_92500_30133# raven_padframe_0|aregc01_3v3_1|GNDR 0.07fF
C9322 raven_padframe_0|aregc01_3v3_1|m4_0_28769# raven_padframe_0|aregc01_3v3_1|GNDO 0.04fF
C9323 raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# 0.17fF
C9324 raven_padframe_0|axtoc02_3v3_0|m4_55000_30653# raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# 0.01fF
C9325 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<12> 1.07fF
C9326 BU_3VX2_63|Q raven_soc_0|gpio_out<11> 0.01fF
C9327 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_outenb<15> 0.02fF
C9328 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<5> 0.01fF
C9329 markings_0|mask_copyright_0|m2_n208_960# markings_0|date_0|_alphabet_2_0|m2_0_0# 0.18fF
C9330 LS_3VX2_19|Q LS_3VX2_22|A 0.16fF
C9331 BU_3VX2_20|A BU_3VX2_19|Q 0.16fF
C9332 BU_3VX2_20|A BU_3VX2_18|Q 0.03fF
C9333 BU_3VX2_73|A vdd 0.05fF
C9334 BU_3VX2_18|A BU_3VX2_15|Q 0.02fF
C9335 LS_3VX2_24|A LS_3VX2_22|A 177.14fF
C9336 raven_soc_0|gpio_pullup<4> BU_3VX2_40|Q 0.22fF
C9337 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<12> 0.02fF
C9338 raven_soc_0|gpio_pullup<7> VDD3V3 0.07fF
C9339 raven_soc_0|gpio_pullup<3> raven_soc_0|ext_clk 0.01fF
C9340 BU_3VX2_0|Q raven_soc_0|gpio_in<8> 0.01fF
C9341 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<11> 20.46fF
C9342 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_in<6> 1.25fF
C9343 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<11> 3.58fF
C9344 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<28> 0.01fF
C9345 BU_3VX2_36|Q BU_3VX2_23|Q 3.50fF
C9346 raven_soc_0|gpio_out<14> apllc03_1v8_0|CLK 0.01fF
C9347 BU_3VX2_71|Q BU_3VX2_23|Q 0.01fF
C9348 BU_3VX2_8|A raven_soc_0|flash_io3_oeb 0.01fF
C9349 BU_3VX2_40|A raven_soc_0|flash_io1_di 0.62fF
C9350 BU_3VX2_17|A BU_3VX2_17|Q 0.08fF
C9351 BU_3VX2_13|A raven_soc_0|flash_io2_do 0.01fF
C9352 raven_soc_0|gpio_out<4> BU_3VX2_71|Q 0.01fF
C9353 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<9> 5.35fF
C9354 raven_soc_0|gpio_in<2> raven_soc_0|flash_io1_di 2.18fF
C9355 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<5> 56.74fF
C9356 LS_3VX2_8|A vdd 3.95fF
C9357 VDD raven_padframe_0|FILLER50F_0|GNDR 0.16fF
C9358 BU_3VX2_0|Q raven_soc_0|gpio_pullup<13> 0.10fF
C9359 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<9> 8.69fF
C9360 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pulldown<7> 3.87fF
C9361 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<8> 0.01fF
C9362 BU_3VX2_27|A raven_soc_0|flash_io1_do 3.71fF
C9363 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<11> 3.93fF
C9364 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<10> 0.02fF
C9365 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<1> 17.40fF
C9366 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<0> 6.55fF
C9367 AMUX2_3V_0|SEL BU_3VX2_49|Q 5.63fF
C9368 BU_3VX2_8|A BU_3VX2_2|A 1.41fF
C9369 BU_3VX2_21|A raven_soc_0|flash_io1_oeb 0.01fF
C9370 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<6> 0.01fF
C9371 raven_padframe_0|BBCUD4F_11|VDDR raven_padframe_0|BBCUD4F_11|GNDR 0.68fF
C9372 raven_soc_0|gpio_in<0> BU_3VX2_27|Q 0.03fF
C9373 raven_soc_0|flash_csb BU_3VX2_27|Q 12.24fF
C9374 raven_soc_0|ram_wdata<5> vdd 0.55fF
C9375 raven_soc_0|irq_pin AMUX4_3V_0|SEL[0] 63.66fF
C9376 raven_soc_0|ram_wdata<0> vdd 0.42fF
C9377 BU_3VX2_52|A BU_3VX2_54|Q 0.04fF
C9378 BU_3VX2_55|Q BU_3VX2_42|Q 0.02fF
C9379 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<8> 0.01fF
C9380 vdd raven_padframe_0|VDDPADF_0|GNDR 0.16fF
C9381 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_outenb<4> 0.43fF
C9382 IN_3VX2_1|A raven_soc_0|gpio_pullup<10> 0.01fF
C9383 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<15> 1.72fF
C9384 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<6> 3.60fF
C9385 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<5> 0.02fF
C9386 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<14> 0.01fF
C9387 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<9> 0.02fF
C9388 BU_3VX2_0|Q raven_soc_0|gpio_out<5> 0.01fF
C9389 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<5> 1.24fF
C9390 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<6> 0.01fF
C9391 raven_soc_0|gpio_out<1> BU_3VX2_24|Q 0.01fF
C9392 LOGIC0_3V_1|Q raven_spi_0|CSB 2.25fF
C9393 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<14> 0.21fF
C9394 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<0> 0.09fF
C9395 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<4> 0.20fF
C9396 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<21> 0.24fF
C9397 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<7> 0.13fF
C9398 BU_3VX2_19|Q BU_3VX2_14|Q 7.76fF
C9399 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<25> 164.03fF
C9400 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<12> 0.21fF
C9401 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<6> 0.01fF
C9402 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<8> 0.19fF
C9403 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<13> 5.53fF
C9404 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<15> 0.22fF
C9405 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<5> 14.44fF
C9406 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<30> 0.01fF
C9407 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<8> 0.02fF
C9408 BU_3VX2_40|Q raven_soc_0|flash_clk 0.13fF
C9409 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<14> 0.01fF
C9410 BU_3VX2_14|Q BU_3VX2_18|Q 14.33fF
C9411 BU_3VX2_70|Q BU_3VX2_5|Q 2.61fF
C9412 BU_3VX2_32|Q BU_3VX2_68|Q 0.56fF
C9413 LS_3VX2_17|A LS_3VX2_16|A 176.65fF
C9414 LS_3VX2_20|A adc0_data<5> 16.23fF
C9415 vdd BU_3VX2_28|Q 1.14fF
C9416 BU_3VX2_43|Q BU_3VX2_45|Q 76.24fF
C9417 LS_3VX2_10|Q LS_3VX2_9|Q 2.67fF
C9418 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<14> 0.01fF
C9419 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<11> 0.01fF
C9420 raven_padframe_0|aregc01_3v3_0|m4_0_0# raven_padframe_0|aregc01_3v3_0|GNDO 1.24fF
C9421 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_out<13> 0.11fF
C9422 raven_padframe_0|BBCUD4F_2|GNDR raven_padframe_0|BBCUD4F_2|VDDO 0.09fF
C9423 AMUX4_3V_1|AIN1 LS_3VX2_15|Q 0.91fF
C9424 BU_3VX2_10|A vdd 0.06fF
C9425 BU_3VX2_4|A raven_soc_0|ext_clk 0.08fF
C9426 analog_out raven_soc_0|irq_pin 3.32fF
C9427 raven_soc_0|gpio_pulldown<12> vdd 0.15fF
C9428 LS_3VX2_4|A vdd 3.84fF
C9429 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<23> 0.01fF
C9430 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<29> 6.69fF
C9431 raven_soc_0|ser_tx BU_3VX2_60|Q 9.83fF
C9432 BU_3VX2_3|A BU_3VX2_2|Q 0.16fF
C9433 LS_3VX2_9|A BU_3VX2_53|Q 18.59fF
C9434 BU_3VX2_35|A VDD3V3 0.31fF
C9435 VDD raven_padframe_0|FILLER01F_1|VDDR 0.71fF
C9436 LS_3VX2_10|A BU_3VX2_62|Q 0.01fF
C9437 AMUX4_3V_4|AOUT raven_soc_0|ext_clk 8.88fF
C9438 BU_3VX2_0|A vdd 0.06fF
C9439 VDD raven_padframe_0|FILLER01F_0|GNDR 0.16fF
C9440 LS_3VX2_24|A BU_3VX2_60|Q 0.02fF
C9441 BU_3VX2_26|A raven_soc_0|flash_io3_di 0.01fF
C9442 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<9> 5.22fF
C9443 raven_soc_0|gpio_pulldown<15> VDD3V3 2.80fF
C9444 BU_3VX2_31|A BU_3VX2_72|Q 0.85fF
C9445 raven_soc_0|gpio_in<2> BU_3VX2_28|Q 0.01fF
C9446 raven_soc_0|gpio_pulldown<1> apllc03_1v8_0|CLK 0.01fF
C9447 BU_3VX2_63|Q raven_soc_0|gpio_in<12> 0.01fF
C9448 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_3|PO 0.04fF
C9449 raven_soc_0|gpio_out<14> raven_soc_0|gpio_outenb<8> 0.74fF
C9450 BU_3VX2_4|Q BU_3VX2_36|Q 3.90fF
C9451 raven_padframe_0|FILLER10F_1|VDDO raven_padframe_0|FILLER10F_1|GNDO 2.28fF
C9452 raven_padframe_0|ICFC_1|VDDO raven_padframe_0|ICFC_1|GNDO 2.28fF
C9453 raven_padframe_0|BBCUD4F_6|GNDR raven_padframe_0|BBCUD4F_6|VDDO 0.09fF
C9454 BU_3VX2_10|A BU_3VX2_40|A 0.45fF
C9455 LS_3VX2_10|A LS_3VX2_5|A 156.98fF
C9456 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<4> 2.97fF
C9457 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<4> 0.52fF
C9458 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<2> 0.01fF
C9459 BU_3VX2_3|A raven_soc_0|flash_clk 0.01fF
C9460 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<12> 0.01fF
C9461 BU_3VX2_15|A raven_soc_0|flash_clk 0.01fF
C9462 raven_padframe_0|BBCUD4F_15|VDDR raven_padframe_0|BBCUD4F_15|VDDO 0.06fF
C9463 raven_soc_0|gpio_in<3> raven_soc_0|flash_io0_oeb 0.06fF
C9464 BU_3VX2_11|A raven_soc_0|flash_io3_di 0.01fF
C9465 raven_soc_0|flash_csb raven_soc_0|flash_io2_oeb 56.23fF
C9466 raven_soc_0|gpio_in<8> raven_soc_0|irq_pin 0.01fF
C9467 BU_3VX2_3|A BU_3VX2_9|A 1.90fF
C9468 VDD raven_padframe_0|BBCUD4F_13|VDDR 0.71fF
C9469 BU_3VX2_9|A BU_3VX2_15|A 2.10fF
C9470 VDD adc_low 0.06fF
C9471 BU_3VX2_0|A BU_3VX2_40|A 0.83fF
C9472 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<10> 0.01fF
C9473 BU_3VX2_6|A raven_soc_0|flash_csb 0.01fF
C9474 raven_soc_0|gpio_in<4> LS_3VX2_3|A 0.01fF
C9475 raven_spi_0|sdo_enb BU_3VX2_33|A 20.40fF
C9476 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<1> 15.02fF
C9477 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<8> 19.41fF
C9478 raven_soc_0|ram_addr<1> raven_soc_0|ram_addr<9> 6.08fF
C9479 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<19> 0.01fF
C9480 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<1> 0.41fF
C9481 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<29> 0.01fF
C9482 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<16> 0.47fF
C9483 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<17> 0.79fF
C9484 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<15> 0.21fF
C9485 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<13> 1.99fF
C9486 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<25> 0.01fF
C9487 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<26> 0.01fF
C9488 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<0> 0.01fF
C9489 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<31> 0.01fF
C9490 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<21> 0.01fF
C9491 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<22> 0.01fF
C9492 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<22> 32.66fF
C9493 BU_3VX2_73|Q LS_3VX2_27|A 57.62fF
C9494 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<16> 0.01fF
C9495 raven_soc_0|ram_wdata<14> raven_soc_0|ram_rdata<13> 0.02fF
C9496 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<29> 38.19fF
C9497 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<1> 0.01fF
C9498 BU_3VX2_51|A BU_3VX2_44|A 0.36fF
C9499 comp_inp vdd 10.09fF
C9500 raven_soc_0|gpio_in<10> BU_3VX2_25|Q 0.01fF
C9501 raven_soc_0|gpio_in<13> BU_3VX2_27|Q 0.01fF
C9502 raven_soc_0|gpio_in<11> BU_3VX2_28|Q 0.01fF
C9503 BU_3VX2_44|Q vdd 1.78fF
C9504 BU_3VX2_45|Q BU_3VX2_50|Q 20.44fF
C9505 raven_padframe_0|BBCUD4F_13|VDDR LOGIC0_3V_4|Q 0.01fF
C9506 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<4> 0.01fF
C9507 raven_padframe_0|aregc01_3v3_1|m4_92500_29333# raven_padframe_0|aregc01_3v3_1|m4_92500_22024# 0.01fF
C9508 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<12> 0.04fF
C9509 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<14> 79.27fF
C9510 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<6> 0.01fF
C9511 LS_3VX2_7|A BU_3VX2_51|Q 0.14fF
C9512 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<11> 14.83fF
C9513 LS_3VX2_3|A raven_soc_0|gpio_in<7> 0.55fF
C9514 BU_3VX2_0|Q VDD3V3 1.86fF
C9515 adc_high BU_3VX2_55|Q 0.13fF
C9516 raven_soc_0|gpio_pulldown<5> raven_soc_0|ext_clk 0.01fF
C9517 raven_soc_0|gpio_out<10> BU_3VX2_29|Q 0.01fF
C9518 raven_soc_0|gpio_pullup<14> BU_3VX2_23|Q 0.01fF
C9519 raven_soc_0|gpio_outenb<9> BU_3VX2_28|Q 0.01fF
C9520 raven_soc_0|gpio_outenb<13> BU_3VX2_26|Q 0.01fF
C9521 BU_3VX2_14|Q BU_3VX2_27|Q 4.98fF
C9522 AMUX4_3V_4|SEL[0] vdd 3.11fF
C9523 BU_3VX2_70|Q BU_3VX2_28|Q 1.20fF
C9524 BU_3VX2_11|Q BU_3VX2_26|Q 0.01fF
C9525 BU_3VX2_7|A raven_soc_0|flash_io0_do 0.01fF
C9526 BU_3VX2_20|A raven_soc_0|flash_io2_oeb 0.01fF
C9527 raven_padframe_0|BT4F_1|VDDR raven_padframe_0|BT4F_1|VDDO 0.06fF
C9528 raven_padframe_0|VDDPADF_1|VDDR raven_padframe_0|VDDPADF_1|GNDR 0.68fF
C9529 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<6> 3.07fF
C9530 raven_soc_0|gpio_pulldown<0> VDD3V3 2.34fF
C9531 raven_spi_0|sdo_enb raven_soc_0|flash_io3_do 0.97fF
C9532 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<14> 0.01fF
C9533 BU_3VX2_33|A raven_soc_0|gpio_in<15> 3.15fF
C9534 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pulldown<7> 6.18fF
C9535 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<12> 0.19fF
C9536 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<9> 0.01fF
C9537 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<19> 132.14fF
C9538 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<23> 3.37fF
C9539 BU_3VX2_49|A BU_3VX2_46|A 1.07fF
C9540 adc0_data<5> BU_3VX2_47|Q 214.90fF
C9541 BU_3VX2_6|A BU_3VX2_20|A 0.01fF
C9542 LS_3VX2_7|Q LS_3VX2_7|A 0.05fF
C9543 BU_3VX2_63|A BU_3VX2_26|A 0.01fF
C9544 BU_3VX2_23|A raven_soc_0|flash_io2_di 0.01fF
C9545 raven_soc_0|gpio_out<0> apllc03_1v8_0|CLK 0.02fF
C9546 raven_padframe_0|ICFC_1|VDDR raven_padframe_0|ICFC_1|VDDO 0.06fF
C9547 BU_3VX2_17|A raven_soc_0|flash_io0_di 0.09fF
C9548 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<6> 0.02fF
C9549 LS_3VX2_13|A LS_3VX2_19|A 0.01fF
C9550 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<6> 0.01fF
C9551 raven_soc_0|gpio_in<0> BU_3VX2_25|Q 0.01fF
C9552 raven_soc_0|ram_wdata<4> vdd 0.52fF
C9553 raven_soc_0|flash_csb BU_3VX2_25|Q 0.01fF
C9554 raven_soc_0|gpio_out<11> BU_3VX2_24|Q 0.01fF
C9555 LS_3VX2_13|A BU_3VX2_52|Q 6.72fF
C9556 raven_soc_0|gpio_out<12> apllc03_1v8_0|CLK 0.01fF
C9557 raven_soc_0|gpio_out<9> BU_3VX2_29|Q 0.01fF
C9558 LOGIC0_3V_1|Q LOGIC1_3V_2|Q 0.21fF
C9559 BU_3VX2_57|A BU_3VX2_57|Q 0.10fF
C9560 BU_3VX2_3|A BU_3VX2_28|A 0.01fF
C9561 BU_3VX2_63|A BU_3VX2_11|A 0.01fF
C9562 BU_3VX2_15|A BU_3VX2_28|A 1.57fF
C9563 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<11> 0.01fF
C9564 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<11> 7.22fF
C9565 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<8> 12.92fF
C9566 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<9> 1.94fF
C9567 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<15> 1.84fF
C9568 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<10> 0.11fF
C9569 LS_3VX2_3|A raven_soc_0|gpio_out<7> 0.01fF
C9570 BU_3VX2_0|Q raven_soc_0|gpio_outenb<6> 0.01fF
C9571 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<10> 0.02fF
C9572 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<14> 0.02fF
C9573 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<6> 11.98fF
C9574 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<31> 0.11fF
C9575 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<6> 0.01fF
C9576 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<7> 0.50fF
C9577 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<0> 0.06fF
C9578 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<12> 4.74fF
C9579 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<24> 0.05fF
C9580 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<2> 0.07fF
C9581 AMUX4_3V_3|SEL[1] BU_3VX2_9|Q 1.38fF
C9582 raven_soc_0|ext_clk raven_soc_0|flash_io0_oeb 39.38fF
C9583 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<5> 0.01fF
C9584 raven_soc_0|flash_io3_di VDD3V3 10.74fF
C9585 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<11> 0.01fF
C9586 raven_padframe_0|aregc01_3v3_0|m4_92500_28769# raven_padframe_0|aregc01_3v3_0|m4_92500_22024# 0.03fF
C9587 raven_padframe_0|aregc01_3v3_0|m4_92500_30653# raven_padframe_0|aregc01_3v3_0|VDDR 0.07fF
C9588 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_outenb<15> 1.11fF
C9589 BU_3VX2_27|A raven_soc_0|flash_csb 9.81fF
C9590 AMUX4_3V_1|AIN1 BU_3VX2_52|A 0.02fF
C9591 AMUX4_3V_4|AIN1 raven_soc_0|irq_pin 2.10fF
C9592 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<2> 3.61fF
C9593 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<21> 0.02fF
C9594 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<15> 20.77fF
C9595 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<0> 0.05fF
C9596 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<25> 0.14fF
C9597 raven_soc_0|ser_tx BU_3VX2_62|Q 18.22fF
C9598 raven_soc_0|ram_rdata<6> vdd 0.16fF
C9599 BU_3VX2_40|A vdd 0.42fF
C9600 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<5> 0.41fF
C9601 LS_3VX2_5|A raven_soc_0|ser_tx 0.01fF
C9602 BU_3VX2_12|A raven_soc_0|flash_io0_di 0.01fF
C9603 LS_3VX2_24|A BU_3VX2_62|Q 0.02fF
C9604 raven_soc_0|ser_rx LS_3VX2_19|A 8.64fF
C9605 IN_3VX2_1|A BU_3VX2_55|Q 0.01fF
C9606 raven_soc_0|gpio_in<2> vdd 3.43fF
C9607 raven_soc_0|gpio_outenb<1> BU_3VX2_27|Q 0.11fF
C9608 raven_soc_0|gpio_out<8> BU_3VX2_71|Q 0.63fF
C9609 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<10> 0.53fF
C9610 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<7> 0.16fF
C9611 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<24> 23.58fF
C9612 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<31> 11.19fF
C9613 BU_3VX2_3|Q BU_3VX2_36|Q 0.10fF
C9614 raven_padframe_0|BBC4F_2|GNDR raven_padframe_0|BBC4F_2|GNDO 0.81fF
C9615 raven_padframe_0|BT4F_0|VDDO raven_padframe_0|BT4F_0|GNDO 2.28fF
C9616 raven_padframe_0|BBCUD4F_8|GNDR raven_padframe_0|BBCUD4F_8|GNDO 0.81fF
C9617 markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# markings_0|manufacturer_0|_alphabet_F_0|m2_0_0# 0.21fF
C9618 BU_3VX2_1|A BU_3VX2_70|A 0.55fF
C9619 LS_3VX2_24|A LS_3VX2_5|A 8.02fF
C9620 raven_soc_0|gpio_pullup<2> BU_3VX2_28|Q 0.01fF
C9621 IN_3VX2_1|A raven_soc_0|flash_io2_di 3.48fF
C9622 raven_soc_0|gpio_in<3> raven_soc_0|flash_io2_do 8.38fF
C9623 raven_soc_0|gpio_out<11> raven_soc_0|gpio_out<15> 0.96fF
C9624 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<7> 0.20fF
C9625 LOGIC0_3V_1|Q BU_3VX2_2|A 0.25fF
C9626 raven_soc_0|irq_pin VDD3V3 7.79fF
C9627 raven_spi_0|SDO LOGIC0_3V_3|Q 1.72fF
C9628 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<12> 0.01fF
C9629 BU_3VX2_20|A BU_3VX2_27|A 3.06fF
C9630 adc_low raven_soc_0|ser_rx 0.05fF
C9631 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<8> 0.01fF
C9632 AMUX4_3V_0|AIN1 BU_3VX2_45|A 0.02fF
C9633 LS_3VX2_12|A BU_3VX2_59|Q 0.01fF
C9634 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<5> 0.92fF
C9635 raven_soc_0|gpio_out<13> raven_soc_0|gpio_out<14> 28.82fF
C9636 raven_soc_0|gpio_out<12> raven_soc_0|gpio_outenb<8> 0.02fF
C9637 raven_soc_0|gpio_out<6> BU_3VX2_71|Q 0.01fF
C9638 LS_3VX2_13|A BU_3VX2_58|Q 0.01fF
C9639 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<1> 14.90fF
C9640 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<5> 5.21fF
C9641 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<8> 0.01fF
C9642 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<9> 0.01fF
C9643 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<6> 3.99fF
C9644 BU_3VX2_66|Q BU_3VX2_21|Q 0.67fF
C9645 raven_soc_0|ram_rdata<12> raven_soc_0|ram_rdata<17> 9.92fF
C9646 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<26> 0.01fF
C9647 BU_3VX2_2|Q BU_3VX2_17|Q 0.24fF
C9648 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<13> 0.05fF
C9649 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<29> 185.25fF
C9650 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<22> 11.22fF
C9651 BU_3VX2_21|Q BU_3VX2_20|Q 60.37fF
C9652 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<21> 14.25fF
C9653 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<27> 0.01fF
C9654 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<1> 0.01fF
C9655 raven_soc_0|gpio_in<11> vdd 1.41fF
C9656 raven_soc_0|gpio_pullup<5> apllc03_1v8_0|CLK 0.09fF
C9657 BU_3VX2_10|Q BU_3VX2_17|Q 4.82fF
C9658 LS_3VX2_16|Q LS_3VX2_17|A 0.20fF
C9659 raven_soc_0|ext_clk BU_3VX2_29|Q 0.01fF
C9660 BU_3VX2_20|Q BU_3VX2_8|Q 2.55fF
C9661 raven_soc_0|gpio_in<12> BU_3VX2_24|Q 0.01fF
C9662 raven_soc_0|gpio_in<13> BU_3VX2_25|Q 0.01fF
C9663 BU_3VX2_62|A vdd 0.07fF
C9664 BU_3VX2_45|Q BU_3VX2_48|Q 32.36fF
C9665 BU_3VX2_3|A BU_3VX2_14|A 0.89fF
C9666 BU_3VX2_5|A BU_3VX2_17|A 0.88fF
C9667 BU_3VX2_15|A BU_3VX2_14|A 38.78fF
C9668 raven_padframe_0|aregc01_3v3_1|m4_92500_31172# raven_padframe_0|aregc01_3v3_1|m4_92500_30653# 0.09fF
C9669 IN_3VX2_1|A raven_soc_0|gpio_pulldown<11> 0.01fF
C9670 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<0> 0.05fF
C9671 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<15> 24.09fF
C9672 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<8> 0.01fF
C9673 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<10> 0.07fF
C9674 BU_3VX2_7|A BU_3VX2_5|Q 0.03fF
C9675 BU_3VX2_63|A VDD3V3 0.20fF
C9676 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<9> 0.44fF
C9677 LS_3VX2_7|A BU_3VX2_49|Q 0.50fF
C9678 LS_3VX2_3|A BU_3VX2_40|Q 22.22fF
C9679 adc_high BU_3VX2_57|Q 0.09fF
C9680 BU_3VX2_1|Q raven_soc_0|flash_io3_oeb 0.53fF
C9681 raven_soc_0|gpio_outenb<9> vdd 0.17fF
C9682 raven_soc_0|gpio_pullup<13> BU_3VX2_26|Q 0.01fF
C9683 BU_3VX2_14|Q BU_3VX2_25|Q 4.11fF
C9684 BU_3VX2_70|Q vdd 1.54fF
C9685 LS_3VX2_21|A BU_3VX2_43|Q 7.32fF
C9686 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<8> 0.01fF
C9687 BU_3VX2_7|A raven_soc_0|flash_io1_di 0.01fF
C9688 BU_3VX2_19|A BU_3VX2_20|Q 0.03fF
C9689 BU_3VX2_16|A BU_3VX2_15|Q 0.16fF
C9690 BU_3VX2_18|A raven_soc_0|flash_io3_do 0.01fF
C9691 IN_3VX2_1|Q AMUX4_3V_0|SEL[1] 4.58fF
C9692 IN_3VX2_1|Q BU_3VX2_51|Q 0.01fF
C9693 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<11> 0.27fF
C9694 LS_3VX2_6|A VDD3V3 0.52fF
C9695 BU_3VX2_0|Q raven_soc_0|ram_wdata<25> 0.02fF
C9696 BU_3VX2_26|A BU_3VX2_26|Q 0.08fF
C9697 BU_3VX2_51|A BU_3VX2_48|A 2.16fF
C9698 BU_3VX2_46|A BU_3VX2_46|Q 0.10fF
C9699 raven_padframe_0|FILLER20F_0|VDDO raven_padframe_0|FILLER20F_0|GNDO 2.28fF
C9700 raven_soc_0|gpio_out<1> raven_soc_0|gpio_in<3> 1.89fF
C9701 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<9> 0.77fF
C9702 raven_soc_0|gpio_in<1> BU_3VX2_27|Q 0.01fF
C9703 BU_3VX2_31|A raven_soc_0|gpio_pullup<14> 0.01fF
C9704 raven_padframe_0|POWERCUTVDD3FC_1|VDDR raven_padframe_0|POWERCUTVDD3FC_1|GNDO 0.13fF
C9705 VDD raven_padframe_0|BBC4F_0|GNDO 0.07fF
C9706 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<8> 0.48fF
C9707 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<10> 1.94fF
C9708 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<7> 0.01fF
C9709 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<9> 0.01fF
C9710 raven_soc_0|gpio_pulldown<2> BU_3VX2_71|Q 0.01fF
C9711 LS_3VX2_13|A LS_3VX2_22|A 32.27fF
C9712 raven_padframe_0|BBCUD4F_8|VDDR raven_padframe_0|BBCUD4F_8|VDDO 0.06fF
C9713 raven_soc_0|ser_rx BU_3VX2_58|Q 2.23fF
C9714 raven_padframe_0|BBCUD4F_4|VDDR raven_padframe_0|BBCUD4F_4|VDDO 0.06fF
C9715 raven_soc_0|gpio_outenb<12> apllc03_1v8_0|CLK 0.01fF
C9716 raven_soc_0|gpio_outenb<10> BU_3VX2_29|Q 0.01fF
C9717 raven_soc_0|gpio_outenb<14> BU_3VX2_28|Q 0.01fF
C9718 AMUX4_3V_3|SEL[0] VDD3V3 0.71fF
C9719 LOGIC1_3V_3|Q LOGIC1_3V_1|Q 0.27fF
C9720 BU_3VX2_23|A BU_3VX2_38|A 0.01fF
C9721 LS_3VX2_10|A LS_3VX2_11|A 54.74fF
C9722 BU_3VX2_5|A BU_3VX2_12|A 1.55fF
C9723 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<11> 11.08fF
C9724 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<3> 4.10fF
C9725 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<4> 0.06fF
C9726 LS_3VX2_3|A raven_soc_0|gpio_outenb<7> 0.01fF
C9727 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<14> 13.78fF
C9728 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<10> 0.02fF
C9729 BU_3VX2_25|A raven_soc_0|flash_io2_di 0.01fF
C9730 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<15> 0.02fF
C9731 BU_3VX2_0|Q raven_soc_0|gpio_pullup<8> 0.01fF
C9732 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<30> 0.02fF
C9733 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<23> 0.01fF
C9734 raven_soc_0|gpio_in<7> raven_soc_0|gpio_in<10> 2.60fF
C9735 AMUX4_3V_3|SEL[1] BU_3VX2_64|Q 0.25fF
C9736 raven_soc_0|gpio_in<12> raven_soc_0|gpio_out<15> 8.95fF
C9737 BU_3VX2_40|Q raven_soc_0|flash_io1_do 0.02fF
C9738 raven_soc_0|ext_clk raven_soc_0|flash_io2_do 21.37fF
C9739 raven_padframe_0|BT4F_2|VDDO raven_padframe_0|BT4F_2|GNDO 2.28fF
C9740 BU_3VX2_0|A BU_3VX2_69|A 0.30fF
C9741 raven_padframe_0|BBCUD4F_5|GNDR raven_padframe_0|BBCUD4F_5|VDDO 0.09fF
C9742 raven_padframe_0|aregc01_3v3_0|m4_92500_31172# raven_padframe_0|aregc01_3v3_0|m4_92500_30133# 0.02fF
C9743 raven_padframe_0|APR00DF_0|VDDO raven_padframe_0|APR00DF_0|GNDO 2.28fF
C9744 BU_3VX2_33|A raven_soc_0|gpio_outenb<15> 4.75fF
C9745 raven_spi_0|SDO VDD3V3 0.17fF
C9746 LS_3VX2_18|Q LS_3VX2_23|Q 46.19fF
C9747 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<28> 58.77fF
C9748 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_pullup<5> 1.04fF
C9749 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<12> 0.27fF
C9750 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<23> 2.13fF
C9751 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<14> 79.43fF
C9752 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<19> 0.26fF
C9753 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<11> 2.48fF
C9754 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<11> 4.90fF
C9755 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<8> 0.01fF
C9756 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<25> 4.45fF
C9757 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<8> 0.01fF
C9758 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<13> 0.01fF
C9759 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<14> 0.01fF
C9760 raven_soc_0|ram_rdata<24> vdd 0.33fF
C9761 BU_3VX2_1|Q apllc03_1v8_0|CLK 2.85fF
C9762 LS_3VX2_21|A BU_3VX2_50|Q 24.43fF
C9763 BU_3VX2_52|Q BU_3VX2_72|Q 1.26fF
C9764 raven_spi_0|CSB LOGIC0_3V_2|Q 1.75fF
C9765 LS_3VX2_12|A AMUX2_3V_0|SEL 23.31fF
C9766 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<0> 8.43fF
C9767 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<14> 0.01fF
C9768 IN_3VX2_1|A BU_3VX2_57|Q 0.01fF
C9769 raven_soc_0|ser_rx LS_3VX2_22|A 0.01fF
C9770 VDD raven_padframe_0|aregc01_3v3_1|m4_0_31172# 0.12fF
C9771 raven_soc_0|gpio_pullup<0> BU_3VX2_23|Q 0.01fF
C9772 BU_3VX2_0|Q BU_3VX2_21|Q 0.01fF
C9773 VDD raven_padframe_0|VDDORPADF_3|GNDO 0.07fF
C9774 VDD raven_padframe_0|APR00DF_2|VDDR 0.71fF
C9775 BU_3VX2_0|Q BU_3VX2_8|Q 0.01fF
C9776 raven_soc_0|gpio_outenb<1> BU_3VX2_25|Q 0.01fF
C9777 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_outenb<13> 43.24fF
C9778 raven_soc_0|gpio_out<8> raven_soc_0|gpio_pullup<14> 0.05fF
C9779 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_out<14> 0.02fF
C9780 raven_soc_0|gpio_pulldown<6> BU_3VX2_71|Q 0.01fF
C9781 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<31> 0.03fF
C9782 raven_soc_0|ram_rdata<30> raven_soc_0|ram_addr<4> 9.63fF
C9783 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<9> 5.35fF
C9784 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<24> 0.18fF
C9785 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<10> 0.41fF
C9786 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<20> 0.88fF
C9787 raven_soc_0|ram_wdata<23> raven_soc_0|ram_addr<2> 0.01fF
C9788 BU_3VX2_10|A BU_3VX2_7|A 5.50fF
C9789 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<15> 1.40fF
C9790 BU_3VX2_3|A raven_soc_0|flash_io1_do 0.01fF
C9791 BU_3VX2_23|A BU_3VX2_23|Q 0.08fF
C9792 raven_soc_0|gpio_pullup<2> vdd 0.35fF
C9793 BU_3VX2_71|A raven_soc_0|flash_io3_do 0.01fF
C9794 BU_3VX2_15|A raven_soc_0|flash_io1_do 0.01fF
C9795 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<7> 0.43fF
C9796 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<15> 1.21fF
C9797 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<10> 1.15fF
C9798 raven_soc_0|gpio_out<11> raven_soc_0|gpio_in<6> 0.33fF
C9799 VDD raven_padframe_0|VDDORPADF_1|GNDO 0.07fF
C9800 BU_3VX2_7|A BU_3VX2_0|A 0.01fF
C9801 BU_3VX2_8|A BU_3VX2_18|A 1.18fF
C9802 LS_3VX2_19|Q acsoc02_3v3_0|CS_4U 0.08fF
C9803 BU_3VX2_38|A IN_3VX2_1|A 0.01fF
C9804 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<2> 8.71fF
C9805 AMUX4_3V_0|AIN1 BU_3VX2_50|A 0.02fF
C9806 LS_3VX2_12|A BU_3VX2_61|Q 0.01fF
C9807 BU_3VX2_11|A BU_3VX2_11|Q 0.08fF
C9808 raven_soc_0|gpio_out<1> raven_soc_0|ext_clk 0.01fF
C9809 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<8> 1.04fF
C9810 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<14> 21.56fF
C9811 raven_soc_0|gpio_out<11> raven_soc_0|gpio_out<10> 17.14fF
C9812 raven_soc_0|gpio_out<5> raven_soc_0|gpio_outenb<13> 0.02fF
C9813 raven_soc_0|gpio_outenb<11> BU_3VX2_71|Q 0.01fF
C9814 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pullup<14> 0.01fF
C9815 LS_3VX2_13|A BU_3VX2_60|Q 0.01fF
C9816 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<27> 1.16fF
C9817 BU_3VX2_15|Q BU_3VX2_38|Q 3.41fF
C9818 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<2> 33.82fF
C9819 BU_3VX2_16|Q BU_3VX2_21|Q 7.00fF
C9820 BU_3VX2_6|Q BU_3VX2_13|Q 8.02fF
C9821 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<29> 1.70fF
C9822 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<25> 6.87fF
C9823 BU_3VX2_19|Q BU_3VX2_66|Q 0.01fF
C9824 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<21> 16.29fF
C9825 raven_soc_0|ram_wdata<14> raven_soc_0|ram_rdata<2> 0.12fF
C9826 BU_3VX2_16|Q BU_3VX2_8|Q 5.10fF
C9827 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<17> 37.48fF
C9828 BU_3VX2_12|Q BU_3VX2_22|Q 5.36fF
C9829 BU_3VX2_21|Q BU_3VX2_30|Q 4.27fF
C9830 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<22> 0.39fF
C9831 BU_3VX2_13|Q BU_3VX2_7|Q 6.93fF
C9832 BU_3VX2_66|Q BU_3VX2_18|Q 0.80fF
C9833 BU_3VX2_19|Q BU_3VX2_20|Q 62.40fF
C9834 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<26> 0.14fF
C9835 BU_3VX2_15|Q BU_3VX2_67|Q 0.04fF
C9836 BU_3VX2_38|Q BU_3VX2_9|Q 3.21fF
C9837 BU_3VX2_73|Q BU_3VX2_53|Q 0.01fF
C9838 BU_3VX2_18|Q BU_3VX2_20|Q 22.17fF
C9839 BU_3VX2_9|Q BU_3VX2_67|Q 7.44fF
C9840 BU_3VX2_55|Q BU_3VX2_54|Q 232.79fF
C9841 BU_3VX2_55|A vdd 0.29fF
C9842 VDD3V3 BU_3VX2_26|Q 1.50fF
C9843 LS_3VX2_21|Q BU_3VX2_44|Q 0.03fF
C9844 LS_3VX2_9|A LS_3VX2_8|A 12.19fF
C9845 raven_padframe_0|FILLER20F_7|VDDR raven_padframe_0|FILLER20F_7|VDDO 0.06fF
C9846 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_in<2> 33.09fF
C9847 BU_3VX2_17|A BU_3VX2_13|A 5.09fF
C9848 raven_padframe_0|aregc01_3v3_1|m4_0_30653# raven_padframe_0|aregc01_3v3_1|m4_0_30133# 0.09fF
C9849 raven_padframe_0|aregc01_3v3_1|m4_0_31172# raven_padframe_0|aregc01_3v3_1|m4_0_29333# 0.01fF
C9850 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<12> 0.02fF
C9851 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<8> 0.75fF
C9852 raven_padframe_0|axtoc02_3v3_0|m4_0_31172# raven_padframe_0|axtoc02_3v3_0|m4_0_30133# 0.03fF
C9853 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<10> 0.01fF
C9854 BU_3VX2_63|Q raven_soc_0|gpio_pullup<4> 0.01fF
C9855 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<3> 0.01fF
C9856 raven_soc_0|ser_tx AMUX4_3V_4|AIN3 45.91fF
C9857 AMUX4_3V_1|SEL[0] BU_3VX2_52|Q 172.92fF
C9858 raven_soc_0|ram_wdata<29> apllc03_1v8_0|CLK 0.01fF
C9859 LS_3VX2_27|A BU_3VX2_43|Q 6.76fF
C9860 LS_3VX2_11|Q LS_3VX2_9|Q 1.16fF
C9861 raven_soc_0|gpio_out<0> raven_soc_0|gpio_out<13> 0.15fF
C9862 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<7> 0.62fF
C9863 raven_soc_0|gpio_in<3> raven_soc_0|gpio_out<11> 0.24fF
C9864 raven_padframe_0|BBCUD4F_1|VDDR raven_padframe_0|BBCUD4F_1|VDDO 0.06fF
C9865 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<8> 0.01fF
C9866 raven_soc_0|gpio_out<12> raven_soc_0|gpio_out<13> 25.48fF
C9867 raven_soc_0|gpio_out<9> raven_soc_0|gpio_out<11> 7.24fF
C9868 BU_3VX2_19|A BU_3VX2_16|Q 0.02fF
C9869 IN_3VX2_1|Q BU_3VX2_49|Q 0.54fF
C9870 BU_3VX2_31|A raven_soc_0|gpio_in<9> 0.01fF
C9871 BU_3VX2_0|Q raven_soc_0|ram_rdata<26> 0.02fF
C9872 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<13> 0.39fF
C9873 LS_3VX2_2|A AMUX4_3V_4|SEL[0] 38.83fF
C9874 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<17> 0.36fF
C9875 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<15> 6.55fF
C9876 raven_soc_0|flash_io0_di raven_soc_0|flash_clk 14.73fF
C9877 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<16> 0.01fF
C9878 BU_3VX2_41|A BU_3VX2_45|Q 0.04fF
C9879 markings_0|date_0|_alphabet_8_0|m2_9_235# markings_0|manufacturer_0|_alphabet_S_1|m2_32_224# 0.17fF
C9880 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<10> 0.03fF
C9881 raven_soc_0|gpio_in<1> BU_3VX2_25|Q 0.01fF
C9882 BU_3VX2_19|A raven_soc_0|flash_io3_di 0.01fF
C9883 BU_3VX2_9|A raven_soc_0|flash_io0_di 0.01fF
C9884 LS_3VX2_11|A raven_soc_0|ser_tx 0.01fF
C9885 BU_3VX2_4|A raven_soc_0|flash_io2_di 0.06fF
C9886 raven_spi_0|SDI raven_padframe_0|ICFC_0|PO 0.04fF
C9887 raven_padframe_0|BT4FC_0|VDD3 raven_padframe_0|BT4FC_0|GNDR 0.16fF
C9888 raven_padframe_0|BT4FC_0|VDDR raven_padframe_0|BT4FC_0|GNDO 0.13fF
C9889 raven_padframe_0|FILLER40F_0|VDDR raven_padframe_0|FILLER40F_0|GNDR 0.68fF
C9890 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<6> 0.21fF
C9891 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<6> 0.03fF
C9892 IN_3VX2_1|A LS_3VX2_16|A 0.01fF
C9893 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<13> 7.35fF
C9894 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<14> 0.41fF
C9895 adc_low AMUX4_3V_1|SEL[0] 0.05fF
C9896 IN_3VX2_1|A BU_3VX2_23|Q 25.95fF
C9897 BU_3VX2_69|A vdd 0.22fF
C9898 raven_soc_0|ser_rx BU_3VX2_60|Q 2.85fF
C9899 raven_soc_0|gpio_outenb<14> vdd 0.21fF
C9900 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_10|PO 0.04fF
C9901 raven_soc_0|gpio_pullup<12> apllc03_1v8_0|CLK 0.01fF
C9902 raven_soc_0|gpio_pullup<15> BU_3VX2_28|Q 0.01fF
C9903 raven_soc_0|gpio_pullup<10> BU_3VX2_29|Q 0.01fF
C9904 LS_3VX2_9|A LS_3VX2_4|A 165.00fF
C9905 LS_3VX2_11|A LS_3VX2_24|A 10.90fF
C9906 BU_3VX2_13|A BU_3VX2_12|A 37.74fF
C9907 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<9> 0.02fF
C9908 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<15> 0.02fF
C9909 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<4> 3.86fF
C9910 LS_3VX2_3|A raven_soc_0|gpio_pullup<9> 0.01fF
C9911 BU_3VX2_63|Q raven_soc_0|flash_clk 0.16fF
C9912 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<7> 0.01fF
C9913 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<15> 0.02fF
C9914 raven_soc_0|gpio_in<12> raven_soc_0|gpio_in<6> 1.11fF
C9915 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<7> 2.82fF
C9916 BU_3VX2_40|Q raven_soc_0|gpio_in<10> 0.06fF
C9917 BU_3VX2_56|A LS_3VX2_17|Q 0.14fF
C9918 BU_3VX2_59|A BU_3VX2_61|A 1.80fF
C9919 BU_3VX2_55|A BU_3VX2_62|A 0.16fF
C9920 BU_3VX2_57|A LS_3VX2_16|Q 0.21fF
C9921 BU_3VX2_58|A LS_3VX2_15|Q 0.35fF
C9922 LS_3VX2_21|Q vdd 0.45fF
C9923 LOGIC0_3V_1|Q raven_spi_0|sdo_enb 3.65fF
C9924 BU_3VX2_8|A BU_3VX2_71|A 0.02fF
C9925 raven_padframe_0|FILLER20FC_0|GNDR raven_padframe_0|FILLER20FC_0|VDDO 0.09fF
C9926 BU_3VX2_38|A BU_3VX2_25|A 0.01fF
C9927 LOGIC1_3V_2|Q LOGIC0_3V_2|Q 0.52fF
C9928 raven_padframe_0|aregc01_3v3_0|m4_0_30653# raven_padframe_0|aregc01_3v3_0|m4_0_29333# 0.02fF
C9929 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<14> 0.01fF
C9930 raven_padframe_0|BBCUD4F_0|GNDR raven_padframe_0|BBCUD4F_0|GNDO 0.81fF
C9931 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<4> 0.01fF
C9932 markings_0|efabless_logo_0|m1_1500_n9450# markings_0|efabless_logo_0|m1_2700_n10050# 0.29fF
C9933 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<9> 5.70fF
C9934 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<20> 0.15fF
C9935 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<11> 0.38fF
C9936 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_out<15> 0.02fF
C9937 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<0> 0.01fF
C9938 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<12> 5.63fF
C9939 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<8> 0.01fF
C9940 LS_3VX2_19|A LS_3VX2_17|A 152.95fF
C9941 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<0> 1.96fF
C9942 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<1> 0.12fF
C9943 raven_soc_0|gpio_outenb<13> VDD3V3 0.07fF
C9944 BU_3VX2_66|Q BU_3VX2_27|Q 3.96fF
C9945 LS_3VX2_2|A vdd 2.77fF
C9946 raven_soc_0|irq_pin adc0_data<5> 11.34fF
C9947 LS_3VX2_27|A BU_3VX2_50|Q 22.23fF
C9948 LS_3VX2_21|A BU_3VX2_48|Q 15.88fF
C9949 LS_3VX2_17|A BU_3VX2_52|Q 7.28fF
C9950 BU_3VX2_20|Q BU_3VX2_27|Q 4.90fF
C9951 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<2> 0.77fF
C9952 BU_3VX2_7|A vdd 0.12fF
C9953 LS_3VX2_14|A BU_3VX2_55|Q 0.02fF
C9954 BU_3VX2_36|A VDD3V3 0.18fF
C9955 BU_3VX2_0|Q BU_3VX2_18|Q 0.01fF
C9956 BU_3VX2_0|Q BU_3VX2_19|Q 0.01fF
C9957 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<4> 4.59fF
C9958 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<30> 0.01fF
C9959 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<8> 2.49fF
C9960 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_pullup<14> 0.02fF
C9961 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<23> 0.01fF
C9962 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<5> 0.05fF
C9963 BU_3VX2_14|Q BU_3VX2_37|Q 2.48fF
C9964 AMUX4_3V_1|SEL[0] BU_3VX2_58|Q 14.10fF
C9965 raven_padframe_0|axtoc02_3v3_0|m4_0_0# raven_padframe_0|axtoc02_3v3_0|GNDO 2.48fF
C9966 BU_3VX2_24|A raven_soc_0|flash_io3_do 0.01fF
C9967 LOGIC0_3V_1|Q raven_soc_0|gpio_in<15> 0.01fF
C9968 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<14> 0.23fF
C9969 BU_3VX2_5|A BU_3VX2_2|Q 0.02fF
C9970 LS_3VX2_10|A LS_3VX2_27|A 5.02fF
C9971 BU_3VX2_67|A BU_3VX2_68|Q 0.03fF
C9972 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<12> 0.04fF
C9973 LS_3VX2_24|A LS_3VX2_21|A 17.97fF
C9974 adc_low LS_3VX2_17|A 0.05fF
C9975 raven_soc_0|gpio_in<0> BU_3VX2_40|Q 0.01fF
C9976 BU_3VX2_28|A raven_soc_0|flash_io0_di 0.01fF
C9977 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<13> 1.23fF
C9978 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<14> 8.91fF
C9979 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<9> 0.36fF
C9980 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<10> 0.25fF
C9981 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<11> 0.11fF
C9982 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<8> 0.27fF
C9983 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<12> 0.03fF
C9984 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<15> 0.48fF
C9985 raven_soc_0|gpio_out<11> raven_soc_0|ext_clk 0.01fF
C9986 raven_soc_0|flash_csb BU_3VX2_40|Q 0.01fF
C9987 raven_soc_0|gpio_out<13> raven_soc_0|gpio_pullup<5> 0.02fF
C9988 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_7|PO 0.04fF
C9989 raven_padframe_0|APR00DF_1|VDDR raven_padframe_0|APR00DF_1|GNDR 0.68fF
C9990 BU_3VX2_7|A BU_3VX2_40|A 0.67fF
C9991 BU_3VX2_19|A BU_3VX2_63|A 0.01fF
C9992 raven_soc_0|gpio_pullup<0> BU_3VX2_31|A 0.01fF
C9993 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<6> 0.01fF
C9994 LS_3VX2_12|A LS_3VX2_15|A 0.16fF
C9995 BU_3VX2_5|A raven_soc_0|flash_clk 0.01fF
C9996 BU_3VX2_25|A BU_3VX2_23|Q 0.03fF
C9997 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_outenb<9> 0.70fF
C9998 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<13> 0.62fF
C9999 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<8> 0.02fF
C10000 BU_3VX2_69|A BU_3VX2_70|Q 0.03fF
C10001 raven_soc_0|gpio_out<5> raven_soc_0|gpio_pullup<13> 0.01fF
C10002 raven_soc_0|gpio_pullup<11> BU_3VX2_71|Q 0.01fF
C10003 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pullup<6> 0.02fF
C10004 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pullup<14> 0.01fF
C10005 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<1> 0.01fF
C10006 raven_soc_0|gpio_pulldown<15> BU_3VX2_27|Q 0.01fF
C10007 LS_3VX2_13|A BU_3VX2_62|Q 0.01fF
C10008 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<14> 36.20fF
C10009 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<3> 0.13fF
C10010 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<12> 0.12fF
C10011 BU_3VX2_16|Q BU_3VX2_19|Q 13.64fF
C10012 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<15> 22.53fF
C10013 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<25> 0.05fF
C10014 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<17> 5.18fF
C10015 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<2> 0.01fF
C10016 BU_3VX2_19|Q BU_3VX2_30|Q 2.49fF
C10017 BU_3VX2_69|Q BU_3VX2_7|Q 0.53fF
C10018 BU_3VX2_38|Q BU_3VX2_64|Q 0.04fF
C10019 BU_3VX2_65|Q BU_3VX2_9|Q 24.96fF
C10020 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<15> 6.33fF
C10021 BU_3VX2_6|Q BU_3VX2_69|Q 1.35fF
C10022 BU_3VX2_30|Q BU_3VX2_18|Q 2.27fF
C10023 BU_3VX2_12|Q BU_3VX2_31|Q 0.02fF
C10024 raven_soc_0|ram_wdata<2> raven_soc_0|ram_wdata<14> 2.02fF
C10025 BU_3VX2_16|Q BU_3VX2_18|Q 22.34fF
C10026 BU_3VX2_68|Q BU_3VX2_10|Q 0.87fF
C10027 BU_3VX2_5|Q BU_3VX2_22|Q 0.98fF
C10028 BU_3VX2_64|Q BU_3VX2_67|Q 4.11fF
C10029 BU_3VX2_2|Q BU_3VX2_68|Q 0.01fF
C10030 VDD3V3 AMUX4_3V_0|SEL[0] 2.31fF
C10031 BU_3VX2_56|Q BU_3VX2_55|Q 230.50fF
C10032 BU_3VX2_57|Q BU_3VX2_54|Q 51.06fF
C10033 LS_3VX2_20|A BU_3VX2_51|Q 158.83fF
C10034 LS_3VX2_20|Q BU_3VX2_43|Q 1.55fF
C10035 AMUX4_3V_0|SEL[1] LS_3VX2_20|A 8.21fF
C10036 raven_padframe_0|CORNERESDF_3|GNDR raven_padframe_0|CORNERESDF_3|VDDO 0.09fF
C10037 BU_3VX2_9|A BU_3VX2_5|A 3.58fF
C10038 LS_3VX2_10|A LS_3VX2_10|Q 0.05fF
C10039 BU_3VX2_23|A BU_3VX2_31|A 4.72fF
C10040 BU_3VX2_2|A LOGIC0_3V_2|Q 0.77fF
C10041 raven_padframe_0|FILLER20F_6|VDDR raven_padframe_0|FILLER20F_6|GNDR 0.68fF
C10042 BU_3VX2_29|A BU_3VX2_33|A 0.02fF
C10043 BU_3VX2_11|A BU_3VX2_26|A 0.01fF
C10044 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<0> 0.21fF
C10045 LS_3VX2_5|A LS_3VX2_13|A 13.41fF
C10046 BU_3VX2_26|A LOGIC0_3V_3|Q 0.19fF
C10047 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<5> 1.23fF
C10048 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<12> 0.01fF
C10049 raven_padframe_0|CORNERESDF_1|GNDR raven_padframe_0|CORNERESDF_1|GNDO 0.81fF
C10050 raven_soc_0|flash_io0_di BU_3VX2_33|Q 0.01fF
C10051 LS_3VX2_22|A AMUX4_3V_1|SEL[0] 0.19fF
C10052 raven_soc_0|ram_wdata<27> vdd 1.30fF
C10053 raven_soc_0|ram_rdata<29> apllc03_1v8_0|CLK 0.01fF
C10054 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<15> 1.36fF
C10055 BU_3VX2_3|A raven_soc_0|flash_csb 0.01fF
C10056 BU_3VX2_15|A raven_soc_0|flash_csb 0.01fF
C10057 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<7> 0.01fF
C10058 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_out<13> 26.49fF
C10059 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_out<11> 18.80fF
C10060 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_out<12> 0.01fF
C10061 analog_out VDD3V3 5.10fF
C10062 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<24> 0.01fF
C10063 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<31> 6.41fF
C10064 raven_soc_0|flash_io3_oeb raven_soc_0|flash_io0_do 351.31fF
C10065 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<17> 3.64fF
C10066 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<16> 15.38fF
C10067 raven_soc_0|flash_io0_oeb raven_soc_0|flash_io2_di 17.05fF
C10068 raven_soc_0|ram_rdata<4> raven_soc_0|ram_addr<0> 0.28fF
C10069 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<22> 57.92fF
C10070 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<27> 4.34fF
C10071 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<25> 0.07fF
C10072 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<15> 86.49fF
C10073 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<13> 0.07fF
C10074 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<31> 0.01fF
C10075 LS_3VX2_17|A BU_3VX2_58|Q 14.41fF
C10076 raven_padframe_0|GNDORPADF_5|VDDO raven_padframe_0|GNDORPADF_5|GNDOR 2.38fF
C10077 raven_padframe_0|FILLER20F_2|GNDR raven_padframe_0|FILLER20F_2|VDDO 0.09fF
C10078 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<10> 0.15fF
C10079 BU_3VX2_2|A raven_soc_0|flash_io0_do 0.01fF
C10080 LS_3VX2_9|A vdd 2.67fF
C10081 BU_3VX2_16|A raven_soc_0|flash_io3_do 0.07fF
C10082 raven_padframe_0|VDDPADFC_0|VDDR raven_padframe_0|VDDPADFC_0|GNDR 0.68fF
C10083 BU_3VX2_29|A raven_soc_0|flash_io3_do 3.77fF
C10084 raven_soc_0|gpio_pullup<8> BU_3VX2_26|Q 0.01fF
C10085 raven_soc_0|gpio_pullup<15> vdd 0.31fF
C10086 raven_soc_0|gpio_outenb<0> apllc03_1v8_0|CLK 0.02fF
C10087 raven_soc_0|ser_rx BU_3VX2_62|Q 4.79fF
C10088 BU_3VX2_0|Q BU_3VX2_27|Q 0.02fF
C10089 BU_3VX2_38|A BU_3VX2_4|A 2.10fF
C10090 LS_3VX2_18|Q LS_3VX2_18|A 0.04fF
C10091 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<3> 12.31fF
C10092 LS_3VX2_5|A raven_soc_0|ser_rx 0.01fF
C10093 BU_3VX2_37|A raven_soc_0|flash_io3_do 0.01fF
C10094 LS_3VX2_3|A raven_soc_0|gpio_pulldown<9> 0.01fF
C10095 BU_3VX2_35|A raven_soc_0|flash_io2_oeb 0.01fF
C10096 LS_3VX2_12|A AMUX4_3V_1|SEL[1] 10.53fF
C10097 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<3> 0.33fF
C10098 BU_3VX2_14|A raven_soc_0|flash_io0_di 0.01fF
C10099 raven_soc_0|gpio_pulldown<0> BU_3VX2_27|Q 0.03fF
C10100 BU_3VX2_24|A BU_3VX2_8|A 0.01fF
C10101 BU_3VX2_40|Q raven_soc_0|gpio_in<13> 0.21fF
C10102 raven_soc_0|ext_clk raven_soc_0|gpio_in<12> 0.01fF
C10103 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<14> 0.02fF
C10104 raven_soc_0|gpio_in<8> VDD3V3 0.07fF
C10105 BU_3VX2_52|A BU_3VX2_58|A 0.69fF
C10106 BU_3VX2_54|A BU_3VX2_56|A 3.67fF
C10107 BU_3VX2_53|A BU_3VX2_57|A 1.23fF
C10108 VDD3V3 BU_3VX2_60|A 0.11fF
C10109 BU_3VX2_3|A BU_3VX2_20|A 0.33fF
C10110 BU_3VX2_6|A BU_3VX2_35|A 0.99fF
C10111 BU_3VX2_20|A BU_3VX2_15|A 3.78fF
C10112 LS_3VX2_12|A LS_3VX2_7|A 153.83fF
C10113 VDD BU_3VX2_33|A 0.02fF
C10114 BU_3VX2_5|A BU_3VX2_28|A 0.01fF
C10115 IN_3VX2_1|A BU_3VX2_31|A 349.69fF
C10116 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<11> 0.02fF
C10117 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<15> 0.01fF
C10118 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<2> 0.01fF
C10119 raven_soc_0|gpio_pulldown<8> BU_3VX2_71|Q 0.01fF
C10120 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<0> 0.01fF
C10121 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_pullup<5> 6.85fF
C10122 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_in<6> 2.53fF
C10123 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<9> 0.02fF
C10124 LS_3VX2_22|A LS_3VX2_17|A 0.01fF
C10125 raven_soc_0|gpio_pullup<13> VDD3V3 0.07fF
C10126 BU_3VX2_6|Q BU_3VX2_29|Q 0.01fF
C10127 BU_3VX2_13|Q BU_3VX2_23|Q 7.13fF
C10128 BU_3VX2_22|Q BU_3VX2_28|Q 6.28fF
C10129 BU_3VX2_2|Q BU_3VX2_24|Q 24.12fF
C10130 BU_3VX2_21|Q BU_3VX2_26|Q 7.84fF
C10131 BU_3VX2_20|Q BU_3VX2_25|Q 7.38fF
C10132 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<4> 2.87fF
C10133 BU_3VX2_10|Q BU_3VX2_24|Q 1.37fF
C10134 BU_3VX2_30|Q BU_3VX2_27|Q 12.32fF
C10135 BU_3VX2_7|Q BU_3VX2_29|Q 1.13fF
C10136 LS_3VX2_16|A BU_3VX2_54|Q 10.99fF
C10137 LS_3VX2_27|Q LS_3VX2_27|A 0.06fF
C10138 BU_3VX2_12|Q apllc03_1v8_0|CLK 0.01fF
C10139 BU_3VX2_8|Q BU_3VX2_26|Q 0.01fF
C10140 BU_3VX2_16|Q BU_3VX2_27|Q 3.17fF
C10141 LS_3VX2_27|A BU_3VX2_48|Q 14.65fF
C10142 BU_3VX2_23|A BU_3VX2_22|A 37.91fF
C10143 LOGIC0_3V_4|Q BU_3VX2_33|A 1.12fF
C10144 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<5> 1.07fF
C10145 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<1> 38.00fF
C10146 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<14> 0.01fF
C10147 LS_3VX2_14|A BU_3VX2_57|Q 0.02fF
C10148 BU_3VX2_26|A VDD3V3 0.58fF
C10149 BU_3VX2_0|Q AMUX4_3V_4|SEL[1] 16.84fF
C10150 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<21> 143.20fF
C10151 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<5> 17.85fF
C10152 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_out<10> 2.99fF
C10153 raven_soc_0|ram_rdata<17> raven_soc_0|ram_rdata<16> 124.78fF
C10154 raven_soc_0|ram_addr<0> raven_soc_0|ram_rdata<15> 2.50fF
C10155 raven_soc_0|ram_rdata<0> vdd 0.36fF
C10156 raven_soc_0|flash_clk BU_3VX2_24|Q 0.01fF
C10157 AMUX4_3V_1|SEL[0] BU_3VX2_60|Q 10.76fF
C10158 raven_soc_0|flash_io3_di BU_3VX2_27|Q 0.01fF
C10159 raven_soc_0|flash_io2_di BU_3VX2_29|Q 0.01fF
C10160 raven_soc_0|flash_io0_do apllc03_1v8_0|CLK 0.01fF
C10161 BU_3VX2_47|Q BU_3VX2_51|Q 34.06fF
C10162 AMUX4_3V_0|SEL[1] BU_3VX2_47|Q 16.20fF
C10163 markings_0|mask_copyright_0|m2_n208_960# markings_0|manufacturer_0|_alphabet_A_1|m2_0_0# 0.14fF
C10164 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<7> 4.43fF
C10165 AMUX4_3V_3|AOUT raven_soc_0|ext_clk 13.42fF
C10166 LS_3VX2_3|Q raven_soc_0|flash_io3_do 0.01fF
C10167 BU_3VX2_13|A BU_3VX2_10|Q 0.02fF
C10168 BU_3VX2_11|A VDD3V3 0.83fF
C10169 raven_padframe_0|ICF_1|VDDR raven_padframe_0|ICF_1|GNDR 0.68fF
C10170 LS_3VX2_24|A LS_3VX2_27|A 25.62fF
C10171 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<15> 8.06fF
C10172 LOGIC0_3V_3|Q VDD3V3 0.38fF
C10173 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<12> 6.53fF
C10174 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<8> 1.03fF
C10175 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<14> 9.40fF
C10176 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<9> 6.75fF
C10177 LS_3VX2_3|A raven_soc_0|flash_io0_di 1.67fF
C10178 BU_3VX2_0|Q raven_soc_0|flash_io2_oeb 0.03fF
C10179 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_pullup<5> 0.02fF
C10180 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<13> 0.02fF
C10181 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<11> 0.01fF
C10182 raven_soc_0|gpio_out<5> VDD3V3 0.07fF
C10183 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<10> 23.31fF
C10184 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<0> 2.80fF
C10185 raven_soc_0|ram_wdata<6> raven_soc_0|ram_rdata<20> 0.38fF
C10186 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<11> 0.05fF
C10187 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<19> 3.47fF
C10188 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<2> 6.97fF
C10189 BU_3VX2_15|A BU_3VX2_14|Q 0.16fF
C10190 IN_3VX2_1|A raven_soc_0|gpio_out<8> 0.01fF
C10191 LOGIC0_3V_4|Q raven_soc_0|flash_io3_do 0.01fF
C10192 BU_3VX2_13|A raven_soc_0|flash_clk 0.01fF
C10193 LOGIC0_3V_4|Q AMUX4_3V_4|AIN3 2.69fF
C10194 raven_soc_0|gpio_out<9> raven_soc_0|gpio_pulldown<7> 5.27fF
C10195 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_pullup<13> 0.24fF
C10196 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<8> 0.15fF
C10197 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<13> 0.10fF
C10198 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pullup<14> 1.50fF
C10199 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<9> 0.02fF
C10200 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<7> 0.01fF
C10201 raven_soc_0|ram_wenb raven_soc_0|ram_addr<6> 0.01fF
C10202 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pullup<6> 0.02fF
C10203 BU_3VX2_33|A raven_soc_0|flash_io1_oeb 0.01fF
C10204 raven_soc_0|gpio_out<3> vdd 0.27fF
C10205 raven_soc_0|gpio_pulldown<14> apllc03_1v8_0|CLK 0.54fF
C10206 raven_soc_0|gpio_pulldown<15> BU_3VX2_25|Q 0.01fF
C10207 raven_soc_0|gpio_pulldown<11> BU_3VX2_29|Q 0.01fF
C10208 raven_padframe_0|BBCUD4F_6|VDDR raven_padframe_0|BBCUD4F_6|VDDO 0.06fF
C10209 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<16> 10.60fF
C10210 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<18> 4.55fF
C10211 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<2> 2.66fF
C10212 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<8> 75.64fF
C10213 BU_3VX2_64|Q BU_3VX2_65|Q 25.76fF
C10214 BU_3VX2_68|Q BU_3VX2_33|Q 0.54fF
C10215 raven_soc_0|ram_wdata<1> raven_soc_0|ram_wdata<8> 3.05fF
C10216 BU_3VX2_57|Q BU_3VX2_56|Q 230.55fF
C10217 BU_3VX2_43|A BU_3VX2_42|Q 0.14fF
C10218 LS_3VX2_20|A BU_3VX2_49|Q 36.01fF
C10219 raven_padframe_0|FILLER40F_0|VDDO raven_padframe_0|FILLER40F_0|GNDO 2.28fF
C10220 BU_3VX2_8|A BU_3VX2_16|A 1.49fF
C10221 raven_padframe_0|CORNERESDF_2|VDDO raven_padframe_0|CORNERESDF_2|GNDO 2.28fF
C10222 BU_3VX2_8|A BU_3VX2_29|A 0.01fF
C10223 BU_3VX2_9|A BU_3VX2_13|A 3.28fF
C10224 raven_padframe_0|VDDORPADF_2|GNDR raven_padframe_0|VDDORPADF_2|GNDO 0.81fF
C10225 LS_3VX2_6|Q LS_3VX2_6|A 0.05fF
C10226 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<10> 0.01fF
C10227 BU_3VX2_63|Q LS_3VX2_3|A 28.43fF
C10228 LOGIC0_3V_4|Q raven_soc_0|gpio_out<14> 9.46fF
C10229 raven_soc_0|ram_addr<1> vdd 0.25fF
C10230 raven_soc_0|ram_wdata<26> vdd 0.85fF
C10231 raven_soc_0|ram_rdata<25> apllc03_1v8_0|CLK 0.01fF
C10232 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<7> 0.15fF
C10233 BU_3VX2_23|A BU_3VX2_21|A 13.14fF
C10234 BU_3VX2_8|A BU_3VX2_37|A 1.11fF
C10235 BU_3VX2_22|A IN_3VX2_1|A 2.68fF
C10236 BU_3VX2_25|A BU_3VX2_31|A 5.64fF
C10237 BU_3VX2_5|A BU_3VX2_14|A 1.19fF
C10238 BU_3VX2_35|A BU_3VX2_27|A 0.01fF
C10239 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<8> 0.13fF
C10240 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<3> 10.40fF
C10241 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<9> 0.01fF
C10242 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_outenb<15> 1.33fF
C10243 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<5> 0.04fF
C10244 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<7> 0.04fF
C10245 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_out<11> 134.94fF
C10246 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_out<13> 182.73fF
C10247 BU_3VX2_73|A BU_3VX2_73|Q 0.10fF
C10248 raven_soc_0|gpio_outenb<1> BU_3VX2_40|Q 0.19fF
C10249 AMUX4_3V_4|AIN1 VDD3V3 2.09fF
C10250 LOGIC0_3V_0|Q raven_spi_0|CSB 2.81fF
C10251 adc_high BU_3VX2_53|A 0.01fF
C10252 raven_soc_0|flash_io3_do raven_soc_0|flash_io1_oeb 34.28fF
C10253 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<13> 5.60fF
C10254 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<10> 0.27fF
C10255 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<17> 15.07fF
C10256 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<13> 0.10fF
C10257 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<1> 5.62fF
C10258 BU_3VX2_13|Q BU_3VX2_4|Q 13.81fF
C10259 BU_3VX2_15|Q BU_3VX2_36|Q 10.21fF
C10260 raven_soc_0|flash_io2_do raven_soc_0|flash_io2_di 81.87fF
C10261 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<24> 0.40fF
C10262 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<29> 3.51fF
C10263 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<7> 0.57fF
C10264 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<2> 0.03fF
C10265 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<21> 150.96fF
C10266 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<26> 2.65fF
C10267 raven_soc_0|flash_io2_oeb raven_soc_0|flash_io3_di 36.86fF
C10268 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<6> 0.08fF
C10269 raven_soc_0|flash_io1_di raven_soc_0|flash_io3_oeb 19.91fF
C10270 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<31> 1.78fF
C10271 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<2> 18.86fF
C10272 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<4> 29.96fF
C10273 raven_soc_0|flash_io1_do raven_soc_0|flash_io0_di 39.93fF
C10274 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<17> 3.04fF
C10275 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<19> 0.01fF
C10276 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<22> 0.01fF
C10277 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<25> 0.01fF
C10278 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<30> 5.66fF
C10279 BU_3VX2_21|Q BU_3VX2_11|Q 3.09fF
C10280 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<27> 0.01fF
C10281 BU_3VX2_36|Q BU_3VX2_9|Q 0.01fF
C10282 BU_3VX2_11|Q BU_3VX2_8|Q 40.69fF
C10283 LS_3VX2_17|A BU_3VX2_60|Q 20.17fF
C10284 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<4> 0.01fF
C10285 BU_3VX2_6|A raven_soc_0|flash_io3_di 0.02fF
C10286 BU_3VX2_2|A raven_soc_0|flash_io1_di 0.02fF
C10287 BU_3VX2_38|A raven_soc_0|flash_io0_oeb 0.01fF
C10288 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<6> 0.23fF
C10289 BU_3VX2_17|A raven_soc_0|ext_clk 0.10fF
C10290 LS_3VX2_14|A LS_3VX2_16|A 0.01fF
C10291 LS_3VX2_8|A BU_3VX2_73|Q 14.53fF
C10292 raven_soc_0|gpio_pulldown<10> apllc03_1v8_0|CLK 0.17fF
C10293 BU_3VX2_0|Q BU_3VX2_25|Q 0.02fF
C10294 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<5> 1.11fF
C10295 BU_3VX2_4|A BU_3VX2_4|Q 0.08fF
C10296 VDD raven_padframe_0|FILLER10F_1|VDDR 0.71fF
C10297 VDD raven_padframe_0|BBCUD4F_14|GNDR 0.16fF
C10298 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<11> 2.65fF
C10299 BU_3VX2_72|A vdd 0.76fF
C10300 BU_3VX2_63|Q raven_soc_0|flash_io1_do 0.03fF
C10301 raven_soc_0|gpio_pulldown<0> BU_3VX2_25|Q 0.01fF
C10302 LS_3VX2_20|Q LS_3VX2_27|Q 4.68fF
C10303 BU_3VX2_43|A BU_3VX2_42|A 1.25fF
C10304 BU_3VX2_8|A LS_3VX2_3|Q 1.28fF
C10305 BU_3VX2_13|A BU_3VX2_28|A 0.01fF
C10306 IN_3VX2_1|A raven_soc_0|gpio_pulldown<2> 0.01fF
C10307 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<7> 0.17fF
C10308 raven_soc_0|gpio_out<2> LS_3VX2_3|A 0.36fF
C10309 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<9> 0.01fF
C10310 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<8> 0.01fF
C10311 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<14> 0.02fF
C10312 raven_soc_0|gpio_pulldown<3> BU_3VX2_40|Q 0.15fF
C10313 raven_soc_0|flash_io2_oeb raven_soc_0|irq_pin 0.01fF
C10314 raven_soc_0|gpio_pulldown<7> raven_soc_0|ext_clk 0.14fF
C10315 BU_3VX2_16|Q BU_3VX2_25|Q 4.00fF
C10316 BU_3VX2_19|Q BU_3VX2_26|Q 7.18fF
C10317 BU_3VX2_35|Q BU_3VX2_29|Q 0.01fF
C10318 BU_3VX2_30|Q BU_3VX2_25|Q 7.61fF
C10319 BU_3VX2_69|Q BU_3VX2_23|Q 12.28fF
C10320 BU_3VX2_22|Q vdd 0.77fF
C10321 BU_3VX2_18|Q BU_3VX2_26|Q 4.37fF
C10322 LS_3VX2_16|A BU_3VX2_56|Q 12.29fF
C10323 BU_3VX2_31|Q BU_3VX2_28|Q 12.26fF
C10324 BU_3VX2_5|Q apllc03_1v8_0|CLK 0.01fF
C10325 VDD3V3 raven_padframe_0|VDDORPADF_4|GNDR 0.78fF
C10326 BU_3VX2_21|A IN_3VX2_1|A 2.33fF
C10327 LS_3VX2_11|A LS_3VX2_13|A 29.84fF
C10328 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<1> 0.01fF
C10329 raven_spi_0|sdo_enb LOGIC0_3V_2|Q 2.58fF
C10330 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<7> 0.01fF
C10331 BU_3VX2_12|A raven_soc_0|ext_clk 0.01fF
C10332 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<16> 0.01fF
C10333 raven_soc_0|ram_rdata<1> raven_soc_0|ram_rdata<13> 1.86fF
C10334 raven_soc_0|ram_wdata<29> raven_soc_0|ram_rdata<15> 0.14fF
C10335 raven_soc_0|ram_wdata<22> raven_soc_0|ram_rdata<16> 0.02fF
C10336 AMUX4_3V_1|SEL[0] BU_3VX2_62|Q 7.93fF
C10337 BU_3VX2_57|A BU_3VX2_58|Q 0.15fF
C10338 BU_3VX2_50|A BU_3VX2_51|Q 0.03fF
C10339 LS_3VX2_15|Q BU_3VX2_59|Q 0.30fF
C10340 raven_soc_0|flash_io3_oeb BU_3VX2_28|Q 0.01fF
C10341 raven_soc_0|flash_io0_oeb BU_3VX2_23|Q 0.01fF
C10342 raven_soc_0|flash_io3_di BU_3VX2_25|Q 0.01fF
C10343 raven_soc_0|flash_io1_di apllc03_1v8_0|CLK 37.20fF
C10344 AMUX4_3V_0|SEL[0] adc0_data<5> 15.43fF
C10345 BU_3VX2_47|Q BU_3VX2_49|Q 74.98fF
C10346 BU_3VX2_45|Q BU_3VX2_72|Q 0.98fF
C10347 BU_3VX2_22|A BU_3VX2_25|A 7.95fF
C10348 raven_padframe_0|BBC4F_3|GNDR raven_padframe_0|BBC4F_3|VDDO 0.09fF
C10349 raven_padframe_0|ICF_0|GNDR raven_padframe_0|ICF_0|GNDO 0.81fF
C10350 raven_padframe_0|FILLER01F_0|VDDO raven_padframe_0|FILLER01F_0|GNDO 2.28fF
C10351 raven_padframe_0|BBCUD4F_9|VDDO raven_padframe_0|BBCUD4F_9|GNDO 2.28fF
C10352 raven_padframe_0|aregc01_3v3_1|m4_0_0# raven_padframe_0|aregc01_3v3_1|GNDO 1.24fF
C10353 raven_padframe_0|axtoc02_3v3_0|m4_0_29057# raven_padframe_0|axtoc02_3v3_0|VDDO 0.07fF
C10354 raven_soc_0|gpio_in<1> BU_3VX2_40|Q 0.01fF
C10355 BU_3VX2_10|A raven_soc_0|flash_io3_oeb 0.01fF
C10356 LS_3VX2_10|A BU_3VX2_53|Q 14.31fF
C10357 BU_3VX2_0|A BU_3VX2_31|Q 0.16fF
C10358 BU_3VX2_20|A BU_3VX2_17|Q 0.02fF
C10359 BU_3VX2_63|A raven_soc_0|flash_io2_oeb 0.01fF
C10360 BU_3VX2_66|A BU_3VX2_66|Q 0.08fF
C10361 VDD raven_padframe_0|APR00DF_5|GNDO 0.07fF
C10362 VDD raven_padframe_0|BBCUD4F_5|GNDR 0.16fF
C10363 LS_3VX2_5|A AMUX4_3V_1|SEL[0] 24.98fF
C10364 raven_soc_0|gpio_outenb<5> BU_3VX2_40|Q 0.82fF
C10365 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<8> 26.59fF
C10366 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<13> 0.02fF
C10367 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<14> 13.35fF
C10368 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<10> 16.61fF
C10369 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<12> 9.75fF
C10370 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<7> 17.81fF
C10371 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<9> 4.77fF
C10372 adc_high BU_3VX2_52|Q 0.45fF
C10373 raven_soc_0|gpio_outenb<6> VDD3V3 0.32fF
C10374 raven_soc_0|ser_rx AMUX4_3V_4|AIN3 64.08fF
C10375 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<20> 0.54fF
C10376 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<19> 27.43fF
C10377 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<0> 0.92fF
C10378 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<23> 60.19fF
C10379 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<11> 0.01fF
C10380 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<28> 6.51fF
C10381 BU_3VX2_10|A BU_3VX2_2|A 0.99fF
C10382 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<11> 0.01fF
C10383 BU_3VX2_6|A BU_3VX2_63|A 0.02fF
C10384 BU_3VX2_8|A raven_soc_0|flash_io1_oeb 0.01fF
C10385 BU_3VX2_5|A raven_soc_0|flash_io1_do 0.01fF
C10386 BU_3VX2_0|A raven_soc_0|flash_io3_oeb 4.54fF
C10387 LS_3VX2_9|Q vdd 1.03fF
C10388 raven_spi_0|sdo_enb raven_soc_0|flash_io0_do 0.63fF
C10389 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<14> 73.46fF
C10390 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<6> 0.70fF
C10391 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<13> 2.57fF
C10392 BU_3VX2_27|A raven_soc_0|flash_io3_di 0.01fF
C10393 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_pulldown<7> 2.99fF
C10394 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<8> 3.78fF
C10395 AMUX4_3V_3|SEL[0] AMUX4_3V_4|SEL[1] 56.28fF
C10396 BU_3VX2_2|A BU_3VX2_0|A 0.03fF
C10397 raven_padframe_0|VDDPADF_0|GNDR raven_padframe_0|VDDPADF_0|VDDO 0.09fF
C10398 BU_3VX2_4|A BU_3VX2_31|A 0.01fF
C10399 LS_3VX2_11|A raven_soc_0|ser_rx 0.01fF
C10400 adc_low adc_high 34.45fF
C10401 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pulldown<12> 0.01fF
C10402 raven_soc_0|gpio_outenb<2> BU_3VX2_71|Q 0.01fF
C10403 LS_3VX2_13|A LS_3VX2_21|A 8.34fF
C10404 LOGIC0_3V_0|Q LOGIC1_3V_2|Q 0.14fF
C10405 BU_3VX2_73|Q comp_inp 1.66fF
C10406 raven_soc_0|ram_wdata<28> vdd 0.74fF
C10407 BU_3VX2_73|Q BU_3VX2_44|Q 7.49fF
C10408 LS_3VX2_22|A BU_3VX2_42|Q 10.88fF
C10409 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<7> 0.01fF
C10410 acsoc02_3v3_0|CS_4U acsoc02_3v3_0|CS_8U 0.32fF
C10411 BU_3VX2_13|A BU_3VX2_14|A 34.78fF
C10412 IN_3VX2_1|A raven_soc_0|gpio_outenb<11> 0.01fF
C10413 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<9> 0.01fF
C10414 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<4> 0.28fF
C10415 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_outenb<15> 9.05fF
C10416 BU_3VX2_0|Q raven_soc_0|ram_wenb 0.25fF
C10417 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<7> 2.09fF
C10418 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<14> 16.83fF
C10419 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_out<13> 0.01fF
C10420 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<7> 7.52fF
C10421 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<5> 0.01fF
C10422 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<8> 1.30fF
C10423 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<3> 7.00fF
C10424 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<10> 0.13fF
C10425 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<4> 0.03fF
C10426 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<20> 0.31fF
C10427 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<31> 0.10fF
C10428 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<6> 3.00fF
C10429 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<24> 5.81fF
C10430 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<18> 0.01fF
C10431 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<2> 0.01fF
C10432 AMUX4_3V_3|SEL[1] BU_3VX2_1|Q 0.97fF
C10433 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<6> 2.76fF
C10434 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<22> 0.01fF
C10435 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<26> 0.01fF
C10436 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<19> 0.03fF
C10437 BU_3VX2_13|Q BU_3VX2_3|Q 12.25fF
C10438 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<2> 0.41fF
C10439 raven_soc_0|ram_wdata<20> raven_soc_0|ram_wdata<14> 10.05fF
C10440 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<21> 0.59fF
C10441 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<22> 0.60fF
C10442 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<8> 24.08fF
C10443 BU_3VX2_6|Q BU_3VX2_32|Q 0.21fF
C10444 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<17> 13.57fF
C10445 BU_3VX2_19|Q BU_3VX2_11|Q 5.46fF
C10446 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<15> 0.01fF
C10447 BU_3VX2_70|Q BU_3VX2_22|Q 25.24fF
C10448 BU_3VX2_32|Q BU_3VX2_7|Q 6.41fF
C10449 BU_3VX2_14|Q BU_3VX2_17|Q 14.47fF
C10450 BU_3VX2_36|Q BU_3VX2_64|Q 17.87fF
C10451 BU_3VX2_4|Q BU_3VX2_69|Q 0.26fF
C10452 BU_3VX2_11|Q BU_3VX2_18|Q 4.77fF
C10453 LS_3VX2_23|A BU_3VX2_33|Q 0.48fF
C10454 LS_3VX2_17|A BU_3VX2_62|Q 59.44fF
C10455 BU_3VX2_26|Q BU_3VX2_27|Q 270.32fF
C10456 BU_3VX2_23|Q BU_3VX2_29|Q 55.62fF
C10457 BU_3VX2_24|Q apllc03_1v8_0|B_CP 0.78fF
C10458 BU_3VX2_28|Q apllc03_1v8_0|CLK 7.49fF
C10459 BU_3VX2_21|A BU_3VX2_25|A 5.60fF
C10460 raven_padframe_0|BBCUD4F_15|GNDR raven_padframe_0|BBCUD4F_15|VDDO 0.09fF
C10461 raven_soc_0|gpio_out<0> LOGIC0_3V_4|Q 0.18fF
C10462 raven_padframe_0|FILLER50F_1|VDDR raven_padframe_0|FILLER50F_1|GNDO 0.13fF
C10463 raven_padframe_0|FILLER50F_1|GNDR raven_padframe_0|FILLER50F_1|VDDO 0.09fF
C10464 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_out<3> 36.20fF
C10465 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pulldown<15> 0.01fF
C10466 LOGIC0_3V_4|Q raven_soc_0|gpio_out<12> 0.01fF
C10467 raven_spi_0|SDO raven_soc_0|flash_io2_oeb 0.42fF
C10468 BU_3VX2_38|A raven_soc_0|flash_io2_do 0.01fF
C10469 LS_3VX2_5|A LS_3VX2_17|A 0.05fF
C10470 VDD raven_padframe_0|BBCUD4F_0|GNDR 0.16fF
C10471 raven_padframe_0|BBCUD4F_5|VDDR raven_padframe_0|BBCUD4F_5|VDDO 0.06fF
C10472 raven_soc_0|gpio_pulldown<12> apllc03_1v8_0|CLK 0.25fF
C10473 LS_3VX2_3|A BU_3VX2_24|Q 0.01fF
C10474 raven_soc_0|ram_rdata<23> raven_soc_0|ram_rdata<17> 12.45fF
C10475 raven_soc_0|ram_rdata<19> raven_soc_0|ram_addr<0> 4.41fF
C10476 AMUX4_3V_0|AIN1 AMUX4_3V_0|SEL[0] 0.02fF
C10477 BU_3VX2_4|A BU_3VX2_3|Q 0.16fF
C10478 IN_3VX2_1|Q BU_3VX2_46|Q 0.88fF
C10479 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<9> 12.77fF
C10480 BU_3VX2_63|Q raven_soc_0|gpio_in<10> 0.07fF
C10481 BU_3VX2_11|A BU_3VX2_8|Q 0.02fF
C10482 IN_3VX2_1|A BU_3VX2_52|Q 0.01fF
C10483 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<15> 35.83fF
C10484 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<7> 0.01fF
C10485 adc_high BU_3VX2_58|Q 0.08fF
C10486 BU_3VX2_0|A BU_3VX2_70|A 0.20fF
C10487 BU_3VX2_19|A BU_3VX2_26|A 3.05fF
C10488 BU_3VX2_63|A BU_3VX2_27|A 0.01fF
C10489 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<13> 0.41fF
C10490 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<3> 4.39fF
C10491 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<9> 0.34fF
C10492 AMUX2_3V_0|AOUT adc_high 2.11fF
C10493 raven_soc_0|gpio_in<0> raven_soc_0|flash_io0_di 0.94fF
C10494 raven_soc_0|gpio_in<3> raven_soc_0|flash_clk 0.11fF
C10495 raven_soc_0|flash_csb raven_soc_0|flash_io0_di 13.55fF
C10496 LOGIC0_3V_0|Q BU_3VX2_2|A 0.38fF
C10497 BU_3VX2_73|Q vdd 7.26fF
C10498 BU_3VX2_31|Q vdd 1.02fF
C10499 AMUX4_3V_4|AIN2 BU_3VX2_55|Q 0.01fF
C10500 BU_3VX2_22|A BU_3VX2_4|A 1.43fF
C10501 BU_3VX2_19|A BU_3VX2_11|A 2.04fF
C10502 IN_3VX2_1|A adc_low 0.05fF
C10503 analog_out LS_3VX2_24|Q 0.02fF
C10504 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<1> 114.99fF
C10505 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<2> 7.23fF
C10506 raven_soc_0|gpio_in<4> BU_3VX2_0|Q 0.01fF
C10507 LOGIC0_3V_1|Q BU_3VX2_37|A 0.03fF
C10508 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<15> 0.12fF
C10509 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<16> 6.08fF
C10510 raven_soc_0|ram_wdata<21> raven_soc_0|ram_rdata<17> 0.02fF
C10511 raven_soc_0|flash_io3_oeb vdd 2.33fF
C10512 raven_soc_0|ext_clk BU_3VX2_59|Q 0.17fF
C10513 BU_3VX2_47|A LS_3VX2_27|Q 0.14fF
C10514 BU_3VX2_46|A BU_3VX2_44|A 2.18fF
C10515 BU_3VX2_41|A LS_3VX2_20|Q 0.27fF
C10516 AMUX4_3V_0|AOUT AMUX4_3V_4|AIN2 1.50fF
C10517 BU_3VX2_57|A BU_3VX2_60|Q 0.02fF
C10518 LS_3VX2_15|Q BU_3VX2_61|Q 1.55fF
C10519 raven_soc_0|flash_io2_do BU_3VX2_23|Q 0.01fF
C10520 raven_soc_0|flash_io1_do BU_3VX2_24|Q 0.01fF
C10521 raven_soc_0|flash_io2_oeb BU_3VX2_26|Q 0.01fF
C10522 BU_3VX2_47|A BU_3VX2_48|Q 0.03fF
C10523 BU_3VX2_50|A BU_3VX2_49|Q 0.15fF
C10524 raven_soc_0|gpio_in<0> BU_3VX2_63|Q 0.01fF
C10525 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<14> 0.41fF
C10526 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<7> 0.01fF
C10527 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_out<11> 31.22fF
C10528 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_out<13> 14.08fF
C10529 BU_3VX2_63|Q raven_soc_0|flash_csb 0.01fF
C10530 BU_3VX2_2|A vdd 0.23fF
C10531 raven_padframe_0|POWERCUTVDD3FC_0|VDDR raven_padframe_0|POWERCUTVDD3FC_0|VDDO 0.06fF
C10532 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<15> 0.02fF
C10533 raven_soc_0|gpio_pullup<7> BU_3VX2_40|Q 0.87fF
C10534 LS_3VX2_24|A BU_3VX2_53|Q 0.01fF
C10535 LS_3VX2_3|A raven_soc_0|gpio_out<15> 0.12fF
C10536 BU_3VX2_0|Q raven_soc_0|gpio_in<7> 0.37fF
C10537 raven_soc_0|gpio_pullup<4> raven_soc_0|ext_clk 0.01fF
C10538 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<13> 0.02fF
C10539 raven_soc_0|gpio_pullup<8> VDD3V3 0.07fF
C10540 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<11> 8.82fF
C10541 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<28> 0.50fF
C10542 raven_padframe_0|FILLER02F_1|VDDR raven_padframe_0|FILLER02F_1|GNDO 0.13fF
C10543 raven_soc_0|gpio_outenb<13> BU_3VX2_27|Q 0.01fF
C10544 raven_soc_0|gpio_outenb<8> BU_3VX2_28|Q 0.01fF
C10545 raven_soc_0|flash_io3_di raven_padframe_0|BBC4F_2|PO 0.04fF
C10546 BU_3VX2_4|Q BU_3VX2_29|Q 0.83fF
C10547 AMUX4_3V_4|SEL[0] apllc03_1v8_0|CLK 17.69fF
C10548 BU_3VX2_11|Q BU_3VX2_27|Q 0.01fF
C10549 BU_3VX2_20|A raven_soc_0|flash_io0_di 0.01fF
C10550 BU_3VX2_40|A raven_soc_0|flash_io3_oeb 0.01fF
C10551 BU_3VX2_18|A raven_soc_0|flash_io0_do 0.01fF
C10552 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<5> 0.01fF
C10553 BU_3VX2_13|A raven_soc_0|flash_io1_do 0.01fF
C10554 raven_spi_0|sdo_enb raven_soc_0|flash_io1_di 2.67fF
C10555 BU_3VX2_31|A raven_soc_0|flash_io0_oeb 42.29fF
C10556 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pulldown<6> 0.15fF
C10557 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<6> 0.37fF
C10558 raven_soc_0|gpio_outenb<4> vdd 0.48fF
C10559 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pulldown<3> 0.01fF
C10560 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<12> 4.03fF
C10561 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<10> 0.06fF
C10562 LS_3VX2_3|A raven_soc_0|gpio_in<5> 0.33fF
C10563 BU_3VX2_0|Q BU_3VX2_37|Q 0.01fF
C10564 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_pulldown<7> 0.02fF
C10565 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<8> 0.69fF
C10566 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<8> 0.01fF
C10567 BU_3VX2_2|A BU_3VX2_40|A 4.11fF
C10568 BU_3VX2_32|A BU_3VX2_36|A 0.51fF
C10569 raven_padframe_0|ICFC_0|VDDR raven_padframe_0|ICFC_0|GNDR 0.68fF
C10570 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<14> 0.42fF
C10571 IN_3VX2_1|A BU_3VX2_58|Q 0.01fF
C10572 LS_3VX2_13|A LS_3VX2_27|A 9.84fF
C10573 raven_soc_0|irq_pin BU_3VX2_51|Q 6.70fF
C10574 BU_3VX2_53|A BU_3VX2_54|Q 0.15fF
C10575 raven_soc_0|irq_pin AMUX4_3V_0|SEL[1] 37.81fF
C10576 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<9> 0.01fF
C10577 BU_3VX2_21|A BU_3VX2_4|A 1.00fF
C10578 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<13> 0.01fF
C10579 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_in<2> 1.14fF
C10580 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<8> 0.01fF
C10581 IN_3VX2_1|A raven_soc_0|gpio_pullup<11> 0.01fF
C10582 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_out<12> 12.32fF
C10583 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<6> 1.77fF
C10584 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_outenb<15> 0.01fF
C10585 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<7> 12.34fF
C10586 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<5> 0.14fF
C10587 BU_3VX2_0|Q raven_soc_0|gpio_out<7> 0.01fF
C10588 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<6> 5.20fF
C10589 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_out<13> 6.43fF
C10590 raven_soc_0|gpio_out<1> BU_3VX2_23|Q 0.01fF
C10591 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<23> 17.45fF
C10592 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<10> 1.13fF
C10593 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<7> 22.50fF
C10594 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<18> 1.17fF
C10595 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<20> 5.24fF
C10596 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<9> 1.06fF
C10597 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<22> 18.04fF
C10598 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<30> 0.22fF
C10599 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<24> 0.01fF
C10600 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<2> 5.75fF
C10601 BU_3VX2_16|Q BU_3VX2_37|Q 4.36fF
C10602 BU_3VX2_3|Q BU_3VX2_69|Q 1.54fF
C10603 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<15> 0.01fF
C10604 raven_soc_0|ram_rdata<21> raven_soc_0|ram_wdata<14> 0.04fF
C10605 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<13> 19.67fF
C10606 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<8> 0.01fF
C10607 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<1> 0.06fF
C10608 raven_soc_0|gpio_out<15> raven_soc_0|flash_io1_do 0.11fF
C10609 BU_3VX2_70|Q BU_3VX2_31|Q 6.29fF
C10610 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<25> 0.01fF
C10611 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<12> 0.18fF
C10612 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<2> 0.04fF
C10613 raven_soc_0|ext_clk raven_soc_0|flash_clk 77.63fF
C10614 raven_soc_0|ram_wdata<7> raven_soc_0|ram_wdata<0> 2.83fF
C10615 VDD3V3 adc0_data<5> 0.02fF
C10616 vdd apllc03_1v8_0|CLK 6.14fF
C10617 BU_3VX2_26|Q BU_3VX2_25|Q 343.12fF
C10618 VDD3V3 raven_padframe_0|VDDORPADF_0|GNDR 0.78fF
C10619 raven_padframe_0|FILLER20FC_0|VDD3 LOGIC0_3V_4|Q 0.04fF
C10620 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<1> 7.29fF
C10621 BU_3VX2_67|A BU_3VX2_65|A 8.42fF
C10622 BU_3VX2_5|A raven_soc_0|flash_csb 0.01fF
C10623 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<4> 2.46fF
C10624 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<12> 0.01fF
C10625 raven_padframe_0|aregc01_3v3_0|m4_92500_0# raven_padframe_0|aregc01_3v3_0|GNDO 1.24fF
C10626 raven_padframe_0|aregc01_3v3_0|VDDR raven_padframe_0|aregc01_3v3_0|GNDR 0.47fF
C10627 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<2> 8.52fF
C10628 BU_3VX2_9|A raven_soc_0|ext_clk 0.01fF
C10629 AMUX4_3V_1|AIN1 LS_3VX2_16|Q 1.07fF
C10630 BU_3VX2_19|A VDD3V3 0.36fF
C10631 VDD raven_padframe_0|BT4F_1|GNDO 0.07fF
C10632 BU_3VX2_70|A vdd 0.25fF
C10633 VDD raven_padframe_0|BBCUD4F_1|GNDO 0.07fF
C10634 BU_3VX2_71|Q raven_soc_0|flash_io3_do 0.32fF
C10635 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<23> 0.01fF
C10636 raven_soc_0|ram_addr<9> raven_soc_0|ram_rdata<19> 0.01fF
C10637 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<13> 0.02fF
C10638 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<27> 3.49fF
C10639 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<29> 0.05fF
C10640 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<31> 0.02fF
C10641 raven_soc_0|ram_rdata<11> raven_soc_0|ram_rdata<1> 1.44fF
C10642 LS_3VX2_21|A BU_3VX2_72|Q 11.48fF
C10643 BU_3VX2_35|A BU_3VX2_40|Q 0.16fF
C10644 LS_3VX2_11|A AMUX4_3V_1|SEL[0] 12.73fF
C10645 LS_3VX2_12|A LS_3VX2_20|A 5.26fF
C10646 VDD raven_padframe_0|BBC4F_3|GNDR 0.16fF
C10647 raven_soc_0|gpio_in<4> raven_soc_0|irq_pin 0.01fF
C10648 raven_soc_0|gpio_pulldown<15> BU_3VX2_40|Q 0.02fF
C10649 BU_3VX2_63|Q raven_soc_0|gpio_in<13> 0.26fF
C10650 BU_3VX2_31|A BU_3VX2_29|Q 63.09fF
C10651 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<14> 221.96fF
C10652 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<12> 24.33fF
C10653 BU_3VX2_27|A BU_3VX2_26|Q 0.16fF
C10654 raven_soc_0|gpio_in<2> apllc03_1v8_0|CLK 0.01fF
C10655 adc_high BU_3VX2_60|Q 0.06fF
C10656 raven_soc_0|gpio_out<14> BU_3VX2_71|Q 0.01fF
C10657 raven_padframe_0|BBCUD4F_6|GNDR raven_padframe_0|BBCUD4F_6|GNDO 0.81fF
C10658 raven_padframe_0|FILLER20F_0|VDDR raven_padframe_0|FILLER20F_0|GNDR 0.68fF
C10659 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<9> 0.01fF
C10660 BU_3VX2_22|A raven_soc_0|flash_io0_oeb 1.76fF
C10661 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<5> 0.48fF
C10662 BU_3VX2_71|A raven_soc_0|flash_io0_do 0.01fF
C10663 raven_padframe_0|BBCUD4F_15|VDDR raven_padframe_0|BBCUD4F_15|GNDO 0.13fF
C10664 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<9> 1.11fF
C10665 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<6> 0.01fF
C10666 raven_padframe_0|FILLER20F_5|VDDR raven_padframe_0|FILLER20F_5|GNDR 0.68fF
C10667 raven_soc_0|gpio_in<7> raven_soc_0|irq_pin 0.01fF
C10668 AMUX4_3V_4|AIN2 BU_3VX2_57|Q 0.01fF
C10669 BU_3VX2_20|A BU_3VX2_5|A 0.01fF
C10670 LOGIC1_3V_3|Q LOGIC0_3V_3|Q 0.52fF
C10671 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<27> 0.03fF
C10672 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<7> 84.05fF
C10673 raven_soc_0|ram_addr<8> raven_soc_0|ram_wdata<21> 0.01fF
C10674 raven_soc_0|ram_rdata<25> raven_soc_0|ram_rdata<15> 5.86fF
C10675 raven_soc_0|ram_wdata<21> raven_soc_0|ram_wdata<22> 156.69fF
C10676 raven_soc_0|ram_wdata<26> raven_soc_0|ram_wdata<27> 174.65fF
C10677 raven_soc_0|ram_rdata<2> raven_soc_0|ram_rdata<1> 39.83fF
C10678 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<31> 0.04fF
C10679 BU_3VX2_1|Q BU_3VX2_67|Q 0.53fF
C10680 raven_soc_0|gpio_in<11> apllc03_1v8_0|CLK 0.02fF
C10681 BU_3VX2_51|A BU_3VX2_43|A 0.25fF
C10682 LS_3VX2_15|Q LS_3VX2_15|A 0.06fF
C10683 raven_soc_0|gpio_in<10> BU_3VX2_24|Q 0.01fF
C10684 LS_3VX2_19|A BU_3VX2_54|Q 7.13fF
C10685 raven_soc_0|gpio_in<15> BU_3VX2_28|Q 0.01fF
C10686 raven_soc_0|gpio_in<8> BU_3VX2_27|Q 0.01fF
C10687 BU_3VX2_54|Q BU_3VX2_52|Q 81.74fF
C10688 BU_3VX2_3|A BU_3VX2_35|A 2.00fF
C10689 raven_padframe_0|aregc01_3v3_1|m4_92500_29057# raven_padframe_0|aregc01_3v3_1|m4_92500_22024# 0.02fF
C10690 raven_padframe_0|aregc01_3v3_1|m4_0_30653# raven_padframe_0|aregc01_3v3_1|VDDR 0.07fF
C10691 IN_3VX2_1|A raven_soc_0|gpio_pulldown<8> 0.01fF
C10692 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<7> 0.01fF
C10693 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_outenb<15> 51.13fF
C10694 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<15> 0.01fF
C10695 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<5> 0.01fF
C10696 BU_3VX2_28|A raven_soc_0|ext_clk 0.01fF
C10697 LS_3VX2_3|A raven_soc_0|gpio_in<6> 0.01fF
C10698 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<15> 0.02fF
C10699 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<14> 0.02fF
C10700 BU_3VX2_0|Q BU_3VX2_40|Q 45.20fF
C10701 BU_3VX2_1|Q raven_soc_0|flash_io1_oeb 0.01fF
C10702 raven_soc_0|gpio_outenb<9> apllc03_1v8_0|CLK 0.01fF
C10703 raven_soc_0|gpio_outenb<8> vdd 0.18fF
C10704 BU_3VX2_11|Q BU_3VX2_25|Q 0.05fF
C10705 raven_soc_0|gpio_outenb<13> BU_3VX2_25|Q 0.01fF
C10706 BU_3VX2_70|Q apllc03_1v8_0|CLK 0.01fF
C10707 raven_soc_0|gpio_out<8> BU_3VX2_29|Q 0.01fF
C10708 BU_3VX2_3|Q BU_3VX2_29|Q 0.01fF
C10709 raven_soc_0|gpio_pullup<13> BU_3VX2_27|Q 0.01fF
C10710 AMUX4_3V_0|AIN1 VDD3V3 3.01fF
C10711 raven_padframe_0|VDDPADF_1|VDDR raven_padframe_0|VDDPADF_1|VDDO 0.06fF
C10712 LS_3VX2_11|A LS_3VX2_17|A 0.01fF
C10713 BU_3VX2_18|A raven_soc_0|flash_io1_di 0.01fF
C10714 raven_padframe_0|BBC4F_2|VDDR raven_padframe_0|BBC4F_2|GNDR 0.68fF
C10715 raven_padframe_0|BT4F_1|VDDR raven_padframe_0|BT4F_1|GNDO 0.13fF
C10716 raven_soc_0|gpio_pulldown<0> BU_3VX2_40|Q 0.33fF
C10717 BU_3VX2_31|A raven_soc_0|flash_io2_do 5.25fF
C10718 BU_3VX2_70|A BU_3VX2_70|Q 0.08fF
C10719 LS_3VX2_8|A BU_3VX2_50|Q 4.65fF
C10720 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pulldown<7> 0.67fF
C10721 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_in<9> 0.02fF
C10722 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pulldown<6> 7.23fF
C10723 LS_3VX2_24|Q VDD3V3 0.69fF
C10724 raven_soc_0|gpio_out<2> raven_soc_0|gpio_in<13> 0.06fF
C10725 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pullup<5> 0.33fF
C10726 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pulldown<3> 1.38fF
C10727 LS_3VX2_3|A raven_soc_0|gpio_out<10> 1.05fF
C10728 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<6> 0.01fF
C10729 adc_low BU_3VX2_54|Q 0.05fF
C10730 BU_3VX2_26|A BU_3VX2_27|Q 0.03fF
C10731 BU_3VX2_47|A BU_3VX2_41|A 9.03fF
C10732 BU_3VX2_48|A BU_3VX2_46|A 1.50fF
C10733 BU_3VX2_49|A BU_3VX2_45|A 0.71fF
C10734 BU_3VX2_49|A BU_3VX2_47|Q 0.04fF
C10735 BU_3VX2_21|A raven_soc_0|flash_io0_oeb 1.59fF
C10736 BU_3VX2_17|A raven_soc_0|flash_io2_di 0.08fF
C10737 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_out<14> 0.01fF
C10738 raven_soc_0|gpio_pulldown<1> BU_3VX2_71|Q 0.20fF
C10739 raven_padframe_0|ICF_0|VDDR raven_padframe_0|ICF_0|VDDO 0.06fF
C10740 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<8> 0.01fF
C10741 IN_3VX2_1|A BU_3VX2_60|Q 0.01fF
C10742 raven_soc_0|gpio_in<0> BU_3VX2_24|Q 0.01fF
C10743 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_9|PO 0.04fF
C10744 raven_soc_0|flash_csb BU_3VX2_24|Q 0.01fF
C10745 raven_soc_0|gpio_out<11> BU_3VX2_23|Q 0.01fF
C10746 raven_soc_0|gpio_out<13> BU_3VX2_28|Q 0.01fF
C10747 raven_soc_0|ext_clk BU_3VX2_33|Q 4.15fF
C10748 raven_soc_0|irq_pin BU_3VX2_49|Q 8.02fF
C10749 BU_3VX2_53|A BU_3VX2_56|Q 0.02fF
C10750 BU_3VX2_58|A BU_3VX2_57|Q 0.03fF
C10751 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<9> 0.01fF
C10752 LS_3VX2_10|A LS_3VX2_8|A 18.13fF
C10753 raven_soc_0|gpio_outenb<1> BU_3VX2_63|Q 0.22fF
C10754 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<9> 6.54fF
C10755 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<10> 0.36fF
C10756 raven_soc_0|gpio_in<3> LS_3VX2_3|A 0.45fF
C10757 LS_3VX2_3|A raven_soc_0|gpio_out<9> 0.01fF
C10758 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_outenb<15> 0.02fF
C10759 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<5> 0.01fF
C10760 BU_3VX2_0|Q raven_soc_0|gpio_outenb<7> 0.01fF
C10761 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<11> 0.02fF
C10762 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<12> 14.77fF
C10763 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_out<13> 64.93fF
C10764 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<10> 0.10fF
C10765 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<7> 12.87fF
C10766 AMUX4_3V_3|SEL[1] BU_3VX2_12|Q 0.05fF
C10767 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<14> 0.36fF
C10768 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<7> 1.50fF
C10769 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<10> 30.58fF
C10770 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<4> 0.05fF
C10771 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<1> 0.10fF
C10772 BU_3VX2_14|Q BU_3VX2_68|Q 18.86fF
C10773 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<2> 0.08fF
C10774 raven_soc_0|gpio_in<10> raven_soc_0|gpio_out<15> 0.65fF
C10775 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<12> 7.67fF
C10776 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<0> 0.01fF
C10777 BU_3VX2_40|Q raven_soc_0|flash_io3_di 11.43fF
C10778 AMUX4_3V_4|AIN2 LS_3VX2_16|A 0.01fF
C10779 BU_3VX2_43|Q BU_3VX2_44|Q 217.86fF
C10780 LS_3VX2_20|A BU_3VX2_46|Q 13.37fF
C10781 BU_3VX2_42|Q BU_3VX2_45|Q 21.62fF
C10782 LOGIC0_3V_0|Q raven_spi_0|sdo_enb 5.25fF
C10783 raven_spi_0|CSB raven_soc_0|gpio_pullup<15> 1.28fF
C10784 VDD3V3 raven_padframe_0|VDDORPADF_1|GNDR 0.78fF
C10785 raven_padframe_0|ICF_1|GNDR raven_padframe_0|ICF_1|GNDO 0.81fF
C10786 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<4> 0.94fF
C10787 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<12> 0.01fF
C10788 raven_padframe_0|aregc01_3v3_0|m4_0_28769# raven_padframe_0|aregc01_3v3_0|GNDO 0.04fF
C10789 BU_3VX2_13|A raven_soc_0|flash_csb 0.01fF
C10790 LOGIC1_3V_3|Q VDD3V3 0.06fF
C10791 AMUX4_3V_1|AIN1 BU_3VX2_53|A 0.02fF
C10792 LS_3VX2_6|Q VDD3V3 0.16fF
C10793 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<23> 31.07fF
C10794 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<10> 0.70fF
C10795 raven_soc_0|ram_rdata<29> raven_soc_0|ram_rdata<19> 7.43fF
C10796 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<0> 0.01fF
C10797 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<11> 0.02fF
C10798 raven_soc_0|ram_addr<7> raven_soc_0|ram_rdata<28> 4.59fF
C10799 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<20> 0.01fF
C10800 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<26> 2.87fF
C10801 raven_soc_0|ram_wdata<7> vdd 0.62fF
C10802 raven_soc_0|ram_rdata<24> apllc03_1v8_0|CLK 0.01fF
C10803 LS_3VX2_27|A BU_3VX2_72|Q 24.18fF
C10804 BU_3VX2_58|Q BU_3VX2_54|Q 34.88fF
C10805 raven_soc_0|gpio_out<1> BU_3VX2_31|A 0.01fF
C10806 LS_3VX2_14|A LS_3VX2_19|A 1.15fF
C10807 LS_3VX2_8|Q VDD3V3 0.16fF
C10808 LS_3VX2_14|A BU_3VX2_52|Q 6.79fF
C10809 BU_3VX2_15|A BU_3VX2_16|Q 0.03fF
C10810 raven_padframe_0|ICFC_0|VDD3 raven_padframe_0|ICFC_0|GNDR 0.16fF
C10811 BU_3VX2_12|A raven_soc_0|flash_io2_di 0.01fF
C10812 BU_3VX2_26|A raven_soc_0|flash_io2_oeb 3.21fF
C10813 BU_3VX2_14|A raven_soc_0|ext_clk 0.01fF
C10814 adc_high BU_3VX2_62|Q 0.05fF
C10815 raven_soc_0|gpio_pulldown<2> BU_3VX2_29|Q 0.01fF
C10816 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_outenb<8> 21.19fF
C10817 raven_soc_0|ram_addr<4> raven_soc_0|ram_rdata<10> 3.09fF
C10818 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<6> 0.11fF
C10819 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<7> 0.18fF
C10820 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<31> 0.14fF
C10821 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<24> 0.01fF
C10822 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_out<14> 33.65fF
C10823 BU_3VX2_32|Q BU_3VX2_4|Q 20.92fF
C10824 raven_soc_0|gpio_in<2> raven_padframe_0|BBCUD4F_2|PO 0.04fF
C10825 raven_padframe_0|FILLER10F_1|VDDR raven_padframe_0|FILLER10F_1|GNDR 0.68fF
C10826 raven_padframe_0|BBCUD4F_14|GNDR raven_padframe_0|BBCUD4F_14|GNDO 0.81fF
C10827 BU_3VX2_10|A BU_3VX2_18|A 1.59fF
C10828 raven_soc_0|gpio_in<1> raven_soc_0|flash_io0_di 0.51fF
C10829 BU_3VX2_24|A raven_soc_0|flash_io0_do 0.01fF
C10830 LOGIC0_3V_0|Q raven_soc_0|gpio_in<15> 0.01fF
C10831 LS_3VX2_10|A LS_3VX2_4|A 33.16fF
C10832 BU_3VX2_6|A BU_3VX2_26|A 0.01fF
C10833 BU_3VX2_3|A raven_soc_0|flash_io3_di 0.01fF
C10834 BU_3VX2_22|A raven_soc_0|flash_io2_do 0.01fF
C10835 raven_soc_0|gpio_pullup<2> apllc03_1v8_0|CLK 0.01fF
C10836 BU_3VX2_71|A raven_soc_0|flash_io1_di 0.01fF
C10837 BU_3VX2_15|A raven_soc_0|flash_io3_di 0.01fF
C10838 BU_3VX2_11|A raven_soc_0|flash_io2_oeb 0.01fF
C10839 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<7> 1.05fF
C10840 raven_soc_0|gpio_in<3> raven_soc_0|flash_io1_do 4.38fF
C10841 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<15> 0.04fF
C10842 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<3> 0.14fF
C10843 VDD raven_padframe_0|BBC4F_0|VDDR 0.71fF
C10844 BU_3VX2_0|A BU_3VX2_18|A 0.01fF
C10845 BU_3VX2_20|A BU_3VX2_13|A 2.45fF
C10846 BU_3VX2_6|A BU_3VX2_11|A 2.31fF
C10847 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_outenb<3> 3.12fF
C10848 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<2> 8.79fF
C10849 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_out<2> 17.41fF
C10850 raven_soc_0|gpio_out<0> BU_3VX2_71|Q 0.12fF
C10851 BU_3VX2_64|A BU_3VX2_36|A 24.48fF
C10852 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<5> 1.31fF
C10853 raven_soc_0|gpio_out<12> BU_3VX2_71|Q 0.01fF
C10854 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<25> 0.02fF
C10855 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<27> 178.72fF
C10856 raven_soc_0|ram_addr<1> raven_soc_0|ram_wdata<26> 0.01fF
C10857 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<1> 0.01fF
C10858 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<22> 1.63fF
C10859 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<17> 0.01fF
C10860 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<31> 5.89fF
C10861 raven_soc_0|ram_wdata<2> raven_soc_0|ram_rdata<1> 0.20fF
C10862 BU_3VX2_20|Q BU_3VX2_17|Q 12.85fF
C10863 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<19> 49.71fF
C10864 LS_3VX2_22|A BU_3VX2_54|Q 0.02fF
C10865 raven_soc_0|ram_wdata<13> raven_soc_0|ram_wdata<25> 4.27fF
C10866 BU_3VX2_66|Q BU_3VX2_17|Q 0.01fF
C10867 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<31> 0.03fF
C10868 BU_3VX2_21|Q BU_3VX2_8|Q 2.30fF
C10869 LS_3VX2_19|A BU_3VX2_56|Q 8.63fF
C10870 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<22> 6.88fF
C10871 BU_3VX2_1|Q BU_3VX2_65|Q 0.51fF
C10872 raven_soc_0|gpio_in<15> vdd 2.01fF
C10873 LS_3VX2_17|Q LS_3VX2_17|A 0.06fF
C10874 raven_soc_0|gpio_in<14> BU_3VX2_28|Q 0.01fF
C10875 raven_soc_0|gpio_in<12> BU_3VX2_23|Q 0.01fF
C10876 raven_soc_0|gpio_in<13> BU_3VX2_24|Q 0.01fF
C10877 BU_3VX2_44|Q BU_3VX2_50|Q 18.36fF
C10878 BU_3VX2_43|Q vdd 1.91fF
C10879 BU_3VX2_56|Q BU_3VX2_52|Q 34.60fF
C10880 raven_soc_0|gpio_in<1> BU_3VX2_63|Q 0.01fF
C10881 VDD3V3 BU_3VX2_27|Q 1.64fF
C10882 LS_3VX2_9|A LS_3VX2_9|Q 0.05fF
C10883 raven_padframe_0|BBC4F_0|VDDR LOGIC0_3V_4|Q 0.01fF
C10884 raven_spi_0|SDI raven_soc_0|gpio_pulldown<15> 1.81fF
C10885 raven_padframe_0|aregc01_3v3_1|m4_92500_31172# raven_padframe_0|aregc01_3v3_1|m4_92500_30133# 0.02fF
C10886 raven_padframe_0|APR00DF_2|VDDO raven_padframe_0|APR00DF_2|GNDO 2.28fF
C10887 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<9> 0.01fF
C10888 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<3> 0.10fF
C10889 raven_padframe_0|axtoc02_3v3_0|m4_0_29333# raven_padframe_0|axtoc02_3v3_0|m4_0_28769# 0.06fF
C10890 BU_3VX2_63|Q raven_soc_0|gpio_outenb<5> 0.01fF
C10891 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<8> 0.33fF
C10892 BU_3VX2_32|A VDD3V3 0.10fF
C10893 BU_3VX2_63|A BU_3VX2_40|Q 0.03fF
C10894 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<12> 0.01fF
C10895 LS_3VX2_3|A raven_soc_0|ext_clk 16.39fF
C10896 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<14> 11.73fF
C10897 raven_soc_0|gpio_pullup<13> BU_3VX2_25|Q 0.01fF
C10898 BU_3VX2_14|Q BU_3VX2_24|Q 5.36fF
C10899 BU_3VX2_37|Q BU_3VX2_26|Q 0.01fF
C10900 BU_3VX2_37|A LOGIC0_3V_2|Q 0.43fF
C10901 BU_3VX2_7|A raven_soc_0|flash_io3_oeb 0.01fF
C10902 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<15> 0.08fF
C10903 adc_low BU_3VX2_56|Q 0.05fF
C10904 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<6> 0.01fF
C10905 raven_padframe_0|BBCUD4F_10|VDDR raven_padframe_0|BBCUD4F_10|VDDO 0.06fF
C10906 BU_3VX2_26|A BU_3VX2_25|Q 0.16fF
C10907 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<11> 3.38fF
C10908 BU_3VX2_50|A BU_3VX2_49|A 12.22fF
C10909 BU_3VX2_45|A BU_3VX2_46|Q 0.03fF
C10910 BU_3VX2_46|Q BU_3VX2_47|Q 76.42fF
C10911 raven_padframe_0|APR00DF_4|VDDR raven_padframe_0|APR00DF_4|GNDR 0.68fF
C10912 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<6> 0.19fF
C10913 BU_3VX2_7|A BU_3VX2_2|A 1.76fF
C10914 BU_3VX2_21|A raven_soc_0|flash_io2_do 0.09fF
C10915 BU_3VX2_16|A raven_soc_0|flash_io0_do 0.05fF
C10916 LS_3VX2_14|A BU_3VX2_58|Q 0.02fF
C10917 BU_3VX2_1|A BU_3VX2_36|Q 0.03fF
C10918 LS_3VX2_8|A raven_soc_0|ser_tx 0.01fF
C10919 raven_padframe_0|ICFC_2|VDD3 raven_padframe_0|ICFC_2|GNDO 0.07fF
C10920 BU_3VX2_13|A BU_3VX2_14|Q 0.03fF
C10921 BU_3VX2_29|A raven_soc_0|flash_io0_do 5.17fF
C10922 IN_3VX2_1|A BU_3VX2_62|Q 0.01fF
C10923 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<3> 1.44fF
C10924 VDD raven_padframe_0|APR00DF_4|VDDR 0.71fF
C10925 raven_soc_0|gpio_outenb<11> BU_3VX2_29|Q 0.01fF
C10926 raven_soc_0|gpio_out<13> vdd 0.23fF
C10927 LS_3VX2_13|A BU_3VX2_53|Q 6.17fF
C10928 raven_soc_0|gpio_outenb<14> apllc03_1v8_0|CLK 0.01fF
C10929 raven_soc_0|gpio_outenb<15> BU_3VX2_28|Q 0.01fF
C10930 AMUX4_3V_4|SEL[1] VDD3V3 0.69fF
C10931 BU_3VX2_3|A BU_3VX2_63|A 0.01fF
C10932 BU_3VX2_10|A BU_3VX2_71|A 0.02fF
C10933 BU_3VX2_63|A BU_3VX2_15|A 0.02fF
C10934 LS_3VX2_2|Q BU_3VX2_1|A 0.01fF
C10935 AMUX4_3V_1|AIN1 adc_low 0.21fF
C10936 LS_3VX2_8|A LS_3VX2_24|A 18.07fF
C10937 BU_3VX2_70|A BU_3VX2_69|A 25.24fF
C10938 BU_3VX2_66|A BU_3VX2_36|A 4.75fF
C10939 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<8> 0.44fF
C10940 BU_3VX2_26|A BU_3VX2_27|A 57.22fF
C10941 BU_3VX2_37|A raven_soc_0|flash_io0_do 0.01fF
C10942 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<12> 30.37fF
C10943 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<4> 6.37fF
C10944 LS_3VX2_3|A raven_soc_0|gpio_outenb<10> 0.01fF
C10945 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<7> 4.87fF
C10946 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_outenb<15> 8.28fF
C10947 BU_3VX2_0|Q raven_soc_0|gpio_pullup<9> 0.01fF
C10948 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<11> 0.02fF
C10949 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<13> 0.01fF
C10950 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<4> 0.27fF
C10951 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<8> 0.07fF
C10952 raven_soc_0|ram_wenb raven_soc_0|ram_addr<3> 0.01fF
C10953 raven_soc_0|gpio_in<11> raven_soc_0|gpio_in<15> 11.18fF
C10954 raven_soc_0|gpio_in<6> raven_soc_0|gpio_in<10> 8.98fF
C10955 raven_soc_0|gpio_in<13> raven_soc_0|gpio_out<15> 16.25fF
C10956 raven_soc_0|ext_clk raven_soc_0|flash_io1_do 21.73fF
C10957 raven_soc_0|flash_io2_oeb VDD3V3 12.02fF
C10958 AMUX4_3V_0|SEL[0] AMUX4_3V_0|SEL[1] 181.66fF
C10959 BU_3VX2_50|Q vdd 2.95fF
C10960 AMUX4_3V_0|SEL[0] BU_3VX2_51|Q 7.97fF
C10961 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<2> 25.56fF
C10962 raven_soc_0|gpio_out<0> raven_soc_0|gpio_outenb<3> 0.38fF
C10963 BU_3VX2_0|A BU_3VX2_71|A 0.01fF
C10964 raven_padframe_0|BBCUD4F_5|GNDR raven_padframe_0|BBCUD4F_5|GNDO 0.81fF
C10965 IN_3VX2_1|A raven_soc_0|gpio_outenb<2> 0.01fF
C10966 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pullup<9> 0.06fF
C10967 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<0> 0.35fF
C10968 BU_3VX2_11|A BU_3VX2_27|A 0.01fF
C10969 BU_3VX2_31|A raven_soc_0|gpio_out<11> 0.01fF
C10970 raven_padframe_0|aregc01_3v3_0|m4_92500_30653# raven_padframe_0|aregc01_3v3_0|m4_92500_30133# 0.09fF
C10971 raven_padframe_0|aregc01_3v3_0|m4_92500_31172# raven_padframe_0|aregc01_3v3_0|m4_92500_29333# 0.01fF
C10972 raven_padframe_0|aregc01_3v3_0|m4_0_29333# raven_padframe_0|aregc01_3v3_0|m4_0_22024# 0.01fF
C10973 raven_soc_0|gpio_in<2> raven_soc_0|gpio_out<13> 0.02fF
C10974 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<5> 0.19fF
C10975 BU_3VX2_6|A VDD3V3 0.30fF
C10976 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<10> 41.56fF
C10977 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<7> 0.04fF
C10978 raven_soc_0|ram_rdata<19> raven_soc_0|ram_rdata<25> 14.37fF
C10979 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<20> 0.65fF
C10980 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<13> 0.93fF
C10981 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<9> 0.53fF
C10982 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<0> 4.56fF
C10983 BU_3VX2_71|Q raven_soc_0|gpio_pullup<5> 0.06fF
C10984 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<15> 0.02fF
C10985 BU_3VX2_59|Q BU_3VX2_55|Q 35.13fF
C10986 raven_soc_0|ram_rdata<4> vdd 0.48fF
C10987 BU_3VX2_1|Q BU_3VX2_72|Q 0.17fF
C10988 BU_3VX2_60|Q BU_3VX2_54|Q 22.00fF
C10989 BU_3VX2_58|Q BU_3VX2_56|Q 82.01fF
C10990 LS_3VX2_2|A apllc03_1v8_0|CLK 1.09fF
C10991 LOGIC0_3V_4|Q LOGIC0_3V_2|Q 0.20fF
C10992 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<2> 6.58fF
C10993 LS_3VX2_9|A BU_3VX2_73|Q 6.72fF
C10994 LS_3VX2_14|A LS_3VX2_22|A 62.61fF
C10995 LS_3VX2_11|A BU_3VX2_42|Q 4.67fF
C10996 LS_3VX2_10|A vdd 2.96fF
C10997 BU_3VX2_18|A vdd 0.06fF
C10998 LS_3VX2_4|A raven_soc_0|ser_tx 0.01fF
C10999 raven_soc_0|gpio_outenb<1> BU_3VX2_24|Q 0.01fF
C11000 BU_3VX2_0|Q BU_3VX2_17|Q 0.01fF
C11001 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<31> 7.90fF
C11002 raven_soc_0|ram_rdata<5> raven_soc_0|ram_rdata<10> 5.87fF
C11003 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<24> 0.60fF
C11004 raven_soc_0|ram_addr<3> raven_soc_0|ram_addr<4> 92.40fF
C11005 raven_soc_0|ram_rdata<30> raven_soc_0|ram_wdata<20> 0.30fF
C11006 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<9> 0.49fF
C11007 raven_soc_0|ram_rdata<8> raven_soc_0|ram_addr<2> 0.65fF
C11008 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<6> 15.84fF
C11009 BU_3VX2_37|Q BU_3VX2_11|Q 21.44fF
C11010 BU_3VX2_3|Q BU_3VX2_32|Q 1.35fF
C11011 raven_padframe_0|APR00DF_1|VDDO raven_padframe_0|APR00DF_1|GNDO 2.28fF
C11012 raven_padframe_0|axtoc02_3v3_0|VDDO raven_padframe_0|axtoc02_3v3_0|GNDO 3.39fF
C11013 markings_0|manufacturer_0|_alphabet_L_0|m2_0_0# markings_0|product_name_0|_alphabet_N_0|m2_0_0# 0.04fF
C11014 BU_3VX2_24|A raven_soc_0|flash_io1_di 0.01fF
C11015 BU_3VX2_38|A BU_3VX2_12|A 1.14fF
C11016 LS_3VX2_24|A LS_3VX2_4|A 6.79fF
C11017 LS_3VX2_3|Q raven_soc_0|flash_io0_do 0.01fF
C11018 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<6> 0.79fF
C11019 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<10> 0.03fF
C11020 IN_3VX2_1|A BU_3VX2_45|Q 9.55fF
C11021 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<10> 8.58fF
C11022 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<11> 11.43fF
C11023 VDD raven_padframe_0|BBCUD4F_5|VDDR 0.71fF
C11024 raven_padframe_0|ICFC_0|VDD3 BU_3VX2_33|A 0.02fF
C11025 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<14> 0.01fF
C11026 LOGIC0_3V_4|Q raven_soc_0|flash_io0_do 0.01fF
C11027 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<10> 0.01fF
C11028 raven_soc_0|gpio_out<12> raven_soc_0|gpio_pullup<14> 0.01fF
C11029 raven_soc_0|gpio_out<11> raven_soc_0|gpio_out<8> 0.85fF
C11030 raven_soc_0|gpio_out<13> raven_soc_0|gpio_outenb<9> 0.21fF
C11031 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_outenb<8> 0.65fF
C11032 raven_soc_0|gpio_outenb<12> BU_3VX2_71|Q 0.01fF
C11033 raven_soc_0|gpio_out<7> raven_soc_0|gpio_outenb<13> 0.01fF
C11034 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<27> 0.70fF
C11035 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<6> 0.01fF
C11036 raven_soc_0|ram_wdata<18> raven_soc_0|ram_addr<5> 0.01fF
C11037 raven_soc_0|ram_wdata<28> raven_soc_0|ram_addr<1> 0.01fF
C11038 BU_3VX2_12|Q BU_3VX2_67|Q 5.69fF
C11039 BU_3VX2_6|Q BU_3VX2_2|Q 11.12fF
C11040 BU_3VX2_19|Q BU_3VX2_21|Q 21.41fF
C11041 BU_3VX2_13|Q BU_3VX2_9|Q 14.15fF
C11042 BU_3VX2_15|Q BU_3VX2_13|Q 22.85fF
C11043 raven_soc_0|ram_rdata<26> raven_soc_0|ram_wdata<13> 0.06fF
C11044 BU_3VX2_19|Q BU_3VX2_8|Q 4.63fF
C11045 BU_3VX2_16|Q BU_3VX2_17|Q 64.14fF
C11046 BU_3VX2_2|Q BU_3VX2_7|Q 8.08fF
C11047 BU_3VX2_6|Q BU_3VX2_10|Q 10.20fF
C11048 BU_3VX2_21|Q BU_3VX2_18|Q 15.50fF
C11049 raven_soc_0|ram_rdata<27> raven_soc_0|ram_wdata<14> 0.01fF
C11050 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<19> 141.85fF
C11051 raven_soc_0|ram_wdata<28> raven_soc_0|ram_wdata<26> 62.87fF
C11052 BU_3VX2_12|Q BU_3VX2_38|Q 2.24fF
C11053 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<17> 5.63fF
C11054 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<25> 3.70fF
C11055 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<19> 3.52fF
C11056 raven_soc_0|ram_wdata<11> raven_soc_0|ram_wdata<22> 4.08fF
C11057 BU_3VX2_18|Q BU_3VX2_8|Q 12.53fF
C11058 BU_3VX2_7|Q BU_3VX2_10|Q 14.22fF
C11059 LS_3VX2_22|A BU_3VX2_56|Q 0.05fF
C11060 BU_3VX2_30|Q BU_3VX2_17|Q 2.05fF
C11061 raven_soc_0|gpio_in<14> vdd 1.45fF
C11062 BU_3VX2_56|A vdd 1.30fF
C11063 BU_3VX2_40|Q BU_3VX2_26|Q 0.01fF
C11064 VDD3V3 BU_3VX2_25|Q 0.79fF
C11065 BU_3VX2_44|Q BU_3VX2_48|Q 25.65fF
C11066 raven_padframe_0|FILLER20F_7|VDDR raven_padframe_0|FILLER20F_7|GNDO 0.13fF
C11067 raven_padframe_0|BBCUD4F_5|VDDR LOGIC0_3V_4|Q 0.01fF
C11068 raven_padframe_0|aregc01_3v3_1|m4_0_30653# raven_padframe_0|aregc01_3v3_1|m4_0_29333# 0.02fF
C11069 raven_padframe_0|APR00DF_2|VDDR raven_padframe_0|APR00DF_2|GNDR 0.68fF
C11070 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<15> 0.39fF
C11071 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<9> 0.70fF
C11072 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<5> 1.30fF
C11073 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<4> 0.01fF
C11074 BU_3VX2_63|Q raven_soc_0|gpio_pullup<7> 0.01fF
C11075 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<6> 0.01fF
C11076 raven_soc_0|gpio_pullup<6> vdd 0.20fF
C11077 AMUX4_3V_3|SEL[1] BU_3VX2_28|Q 0.30fF
C11078 raven_soc_0|ser_tx comp_inp 27.74fF
C11079 raven_soc_0|ram_rdata<15> vdd 0.34fF
C11080 LS_3VX2_21|A BU_3VX2_42|Q 165.72fF
C11081 raven_soc_0|ram_wdata<27> apllc03_1v8_0|CLK 0.01fF
C11082 raven_soc_0|gpio_in<0> raven_soc_0|gpio_in<3> 0.59fF
C11083 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<14> 14.47fF
C11084 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<9> 1.74fF
C11085 raven_padframe_0|BBCUD4F_1|VDDR raven_padframe_0|BBCUD4F_1|GNDO 0.13fF
C11086 raven_soc_0|gpio_out<6> raven_soc_0|gpio_out<11> 0.48fF
C11087 markings_0|product_name_0|_alphabet_E_0|m2_0_0# markings_0|product_name_0|_alphabet_V_0|m2_0_560# 1.23fF
C11088 markings_0|efabless_logo_0|m1_6600_n2850# markings_0|efabless_logo_0|m1_7500_n3450# 0.21fF
C11089 BU_3VX2_19|A BU_3VX2_19|Q 0.08fF
C11090 BU_3VX2_9|A BU_3VX2_6|Q 0.02fF
C11091 BU_3VX2_9|A BU_3VX2_7|Q 0.03fF
C11092 BU_3VX2_19|A BU_3VX2_18|Q 0.16fF
C11093 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<5> 0.24fF
C11094 LS_3VX2_14|Q VDD3V3 0.20fF
C11095 VDD raven_padframe_0|FILLER20F_6|VDDR 0.71fF
C11096 raven_soc_0|gpio_in<2> raven_soc_0|gpio_in<14> 0.41fF
C11097 BU_3VX2_31|A raven_soc_0|gpio_in<12> 0.01fF
C11098 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pulldown<7> 0.01fF
C11099 BU_3VX2_27|A VDD3V3 1.46fF
C11100 adc_high AMUX4_3V_4|AIN3 4.65fF
C11101 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<16> 0.34fF
C11102 raven_soc_0|flash_io0_do raven_soc_0|flash_io1_oeb 91.32fF
C11103 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<13> 16.71fF
C11104 raven_soc_0|ram_rdata<31> raven_soc_0|ram_rdata<17> 0.17fF
C11105 BU_3VX2_1|Q BU_3VX2_36|Q 1.02fF
C11106 raven_soc_0|flash_io2_di raven_soc_0|flash_clk 14.95fF
C11107 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<15> 2.98fF
C11108 raven_padframe_0|BBC4F_0|GNDR raven_padframe_0|BBC4F_0|GNDO 0.81fF
C11109 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<11> 0.18fF
C11110 raven_soc_0|gpio_in<1> BU_3VX2_24|Q 0.01fF
C11111 BU_3VX2_23|A raven_soc_0|flash_io3_do 0.01fF
C11112 BU_3VX2_9|A raven_soc_0|flash_io2_di 0.01fF
C11113 BU_3VX2_16|A raven_soc_0|flash_io1_di 0.09fF
C11114 raven_padframe_0|FILLER40F_0|VDDR raven_padframe_0|FILLER40F_0|VDDO 0.06fF
C11115 LS_3VX2_14|A BU_3VX2_60|Q 0.02fF
C11116 BU_3VX2_71|A vdd 0.13fF
C11117 raven_soc_0|gpio_in<4> raven_soc_0|gpio_in<8> 0.99fF
C11118 BU_3VX2_29|A raven_soc_0|flash_io1_di 0.01fF
C11119 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<6> 0.01fF
C11120 IN_3VX2_1|A apllc03_1v8_0|B_VCO 0.43fF
C11121 VDD raven_padframe_0|FILLER20F_2|GNDR 0.16fF
C11122 raven_padframe_0|BBCUD4F_12|VDDR raven_padframe_0|BBCUD4F_12|GNDR 0.68fF
C11123 AMUX2_3V_0|SEL BU_3VX2_55|Q 0.01fF
C11124 raven_soc_0|gpio_outenb<15> vdd 0.30fF
C11125 raven_soc_0|gpio_pullup<8> BU_3VX2_27|Q 0.01fF
C11126 raven_soc_0|gpio_pullup<11> BU_3VX2_29|Q 0.01fF
C11127 raven_soc_0|gpio_pullup<15> apllc03_1v8_0|CLK 0.01fF
C11128 BU_3VX2_24|A BU_3VX2_10|A 0.01fF
C11129 BU_3VX2_68|A BU_3VX2_33|A 1.21fF
C11130 BU_3VX2_37|A raven_soc_0|flash_io1_di 0.01fF
C11131 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<0> 0.01fF
C11132 LS_3VX2_3|A raven_soc_0|gpio_pullup<10> 0.01fF
C11133 BU_3VX2_35|A raven_soc_0|flash_io0_di 0.14fF
C11134 BU_3VX2_0|Q raven_soc_0|gpio_pulldown<9> 0.01fF
C11135 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<13> 0.01fF
C11136 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<22> 0.04fF
C11137 LOGIC0_3V_4|Q raven_padframe_0|BBC4F_0|PO 0.04fF
C11138 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<10> 4.17fF
C11139 raven_soc_0|gpio_in<13> raven_soc_0|gpio_in<6> 7.04fF
C11140 raven_soc_0|gpio_in<8> raven_soc_0|gpio_in<7> 23.64fF
C11141 raven_soc_0|gpio_in<14> raven_soc_0|gpio_in<11> 1.69fF
C11142 raven_soc_0|ext_clk raven_soc_0|gpio_in<10> 0.01fF
C11143 BU_3VX2_24|A BU_3VX2_0|A 0.01fF
C11144 BU_3VX2_59|A LS_3VX2_15|Q 0.49fF
C11145 BU_3VX2_60|A BU_3VX2_61|A 4.81fF
C11146 BU_3VX2_57|A LS_3VX2_17|Q 0.16fF
C11147 BU_3VX2_56|A BU_3VX2_62|A 0.18fF
C11148 BU_3VX2_58|A LS_3VX2_16|Q 0.25fF
C11149 LS_3VX2_27|Q vdd 0.04fF
C11150 AMUX4_3V_0|SEL[0] BU_3VX2_49|Q 9.89fF
C11151 BU_3VX2_48|Q vdd 2.66fF
C11152 raven_padframe_0|APR00DF_5|VDDR raven_padframe_0|APR00DF_5|VDDO 0.06fF
C11153 BU_3VX2_71|A BU_3VX2_40|A 0.07fF
C11154 raven_padframe_0|BBCUD4F_13|GNDR raven_padframe_0|BBCUD4F_13|GNDO 0.81fF
C11155 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_pulldown<9> 0.28fF
C11156 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<10> 0.01fF
C11157 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<7> 0.01fF
C11158 raven_padframe_0|aregc01_3v3_0|m4_0_30133# raven_padframe_0|aregc01_3v3_0|m4_0_29333# 0.09fF
C11159 raven_padframe_0|aregc01_3v3_0|m4_0_30653# raven_padframe_0|aregc01_3v3_0|m4_0_29057# 0.01fF
C11160 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pullup<3> 1.75fF
C11161 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_outenb<0> 8.28fF
C11162 raven_soc_0|gpio_in<2> raven_soc_0|gpio_outenb<15> 0.01fF
C11163 raven_padframe_0|BBCUD4F_0|VDDO raven_padframe_0|BBCUD4F_0|GNDO 2.28fF
C11164 raven_soc_0|gpio_out<10> raven_soc_0|gpio_in<13> 0.75fF
C11165 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_in<14> 0.03fF
C11166 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<12> 5.80fF
C11167 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_pullup<5> 0.17fF
C11168 raven_soc_0|gpio_outenb<13> BU_3VX2_40|Q 0.31fF
C11169 raven_soc_0|ram_rdata<28> raven_soc_0|ram_wdata<2> 0.01fF
C11170 raven_soc_0|ram_wdata<5> raven_soc_0|ram_rdata<19> 0.20fF
C11171 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<12> 0.24fF
C11172 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<0> 0.39fF
C11173 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_in<11> 0.02fF
C11174 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<7> 0.01fF
C11175 raven_soc_0|ser_tx vdd 4.39fF
C11176 BU_3VX2_21|Q BU_3VX2_27|Q 7.19fF
C11177 BU_3VX2_59|Q BU_3VX2_57|Q 84.86fF
C11178 BU_3VX2_61|Q BU_3VX2_55|Q 22.28fF
C11179 BU_3VX2_62|Q BU_3VX2_54|Q 15.42fF
C11180 BU_3VX2_8|Q BU_3VX2_27|Q 7.44fF
C11181 BU_3VX2_60|Q BU_3VX2_56|Q 34.86fF
C11182 BU_3VX2_53|Q BU_3VX2_72|Q 1.54fF
C11183 BU_3VX2_35|A BU_3VX2_63|Q 0.03fF
C11184 raven_soc_0|gpio_in<4> raven_soc_0|gpio_out<5> 0.15fF
C11185 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_out<3> 1.75fF
C11186 BU_3VX2_63|Q raven_soc_0|gpio_pulldown<15> 0.01fF
C11187 LS_3VX2_19|Q vdd 0.06fF
C11188 LS_3VX2_24|A vdd 4.26fF
C11189 BU_3VX2_64|A VDD3V3 0.07fF
C11190 VDD raven_padframe_0|VDDORPADF_2|GNDR 0.16fF
C11191 LS_3VX2_5|A BU_3VX2_54|Q 13.00fF
C11192 VDD raven_padframe_0|FILLER02F_0|GNDO 0.07fF
C11193 VDD raven_padframe_0|APR00DF_3|GNDO 0.07fF
C11194 VDD raven_padframe_0|CORNERESDF_1|VDDR 0.71fF
C11195 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_outenb<9> 2.31fF
C11196 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<8> 3.49fF
C11197 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<4> 0.32fF
C11198 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<20> 0.14fF
C11199 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<30> 8.94fF
C11200 raven_soc_0|ram_rdata<5> raven_soc_0|ram_addr<3> 0.31fF
C11201 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<23> 0.11fF
C11202 raven_soc_0|ram_rdata<22> raven_soc_0|ram_addr<2> 4.42fF
C11203 AMUX4_3V_3|SEL[1] AMUX4_3V_4|SEL[0] 59.17fF
C11204 raven_padframe_0|ICFC_2|GNDR raven_padframe_0|ICFC_2|VDDO 0.09fF
C11205 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<15> 0.83fF
C11206 raven_soc_0|gpio_out<0> raven_soc_0|gpio_in<9> 0.01fF
C11207 LS_3VX2_3|Q raven_soc_0|flash_io1_di 0.01fF
C11208 IN_3VX2_1|A raven_soc_0|flash_io3_do 4.18fF
C11209 IN_3VX2_1|A AMUX4_3V_4|AIN3 5.16fF
C11210 BU_3VX2_28|A raven_soc_0|flash_io2_di 0.01fF
C11211 raven_soc_0|gpio_in<0> raven_soc_0|ext_clk 0.01fF
C11212 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<10> 116.70fF
C11213 raven_soc_0|gpio_out<7> raven_soc_0|gpio_in<8> 3.69fF
C11214 VDD raven_padframe_0|BBCUD4F_12|GNDO 0.07fF
C11215 raven_soc_0|gpio_out<9> raven_soc_0|gpio_in<13> 0.83fF
C11216 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<15> 21.76fF
C11217 raven_soc_0|gpio_out<5> raven_soc_0|gpio_in<7> 1.74fF
C11218 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_in<11> 0.21fF
C11219 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<12> 0.03fF
C11220 raven_soc_0|gpio_out<12> raven_soc_0|gpio_in<9> 7.33fF
C11221 BU_3VX2_0|Q raven_soc_0|flash_io0_di 14.58fF
C11222 BU_3VX2_29|A BU_3VX2_28|Q 0.16fF
C11223 raven_soc_0|flash_csb raven_soc_0|ext_clk 176.01fF
C11224 raven_soc_0|gpio_in<3> raven_soc_0|gpio_in<13> 0.01fF
C11225 raven_spi_0|SDO raven_spi_0|SDI 24.04fF
C11226 BU_3VX2_10|A BU_3VX2_16|A 2.16fF
C11227 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<5> 5.42fF
C11228 BU_3VX2_10|A BU_3VX2_29|A 0.01fF
C11229 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<1> 18.54fF
C11230 LOGIC0_3V_4|Q raven_soc_0|flash_io1_di 0.10fF
C11231 IN_3VX2_1|A raven_soc_0|gpio_out<14> 0.01fF
C11232 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<8> 0.02fF
C11233 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_outenb<13> 0.76fF
C11234 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_outenb<9> 0.54fF
C11235 raven_soc_0|gpio_pullup<12> BU_3VX2_71|Q 0.01fF
C11236 raven_soc_0|gpio_out<7> raven_soc_0|gpio_pullup<13> 0.01fF
C11237 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_pullup<14> 7.71fF
C11238 raven_soc_0|gpio_out<11> raven_soc_0|gpio_pulldown<6> 0.02fF
C11239 raven_padframe_0|BBCUD4F_9|VDDR raven_padframe_0|BBCUD4F_9|GNDO 0.13fF
C11240 raven_soc_0|gpio_out<3> apllc03_1v8_0|CLK 0.01fF
C11241 raven_soc_0|gpio_pulldown<8> BU_3VX2_29|Q 0.01fF
C11242 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<30> 6.41fF
C11243 raven_soc_0|ram_wdata<11> raven_soc_0|ram_rdata<27> 0.31fF
C11244 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<26> 0.45fF
C11245 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<29> 0.49fF
C11246 BU_3VX2_38|Q BU_3VX2_5|Q 13.32fF
C11247 BU_3VX2_19|Q BU_3VX2_18|Q 67.36fF
C11248 BU_3VX2_12|Q BU_3VX2_65|Q 2.15fF
C11249 BU_3VX2_15|Q BU_3VX2_69|Q 0.16fF
C11250 BU_3VX2_13|Q BU_3VX2_64|Q 0.19fF
C11251 BU_3VX2_66|Q BU_3VX2_68|Q 8.12fF
C11252 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<15> 0.27fF
C11253 raven_soc_0|ram_wdata<12> raven_soc_0|ram_wdata<13> 92.79fF
C11254 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<17> 0.26fF
C11255 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<1> 0.01fF
C11256 BU_3VX2_35|Q BU_3VX2_2|Q 10.76fF
C11257 BU_3VX2_35|Q BU_3VX2_10|Q 2.17fF
C11258 BU_3VX2_69|Q BU_3VX2_9|Q 2.24fF
C11259 BU_3VX2_68|Q BU_3VX2_20|Q 0.01fF
C11260 BU_3VX2_31|Q BU_3VX2_22|Q 3.37fF
C11261 BU_3VX2_33|Q BU_3VX2_7|Q 0.01fF
C11262 BU_3VX2_5|Q BU_3VX2_67|Q 0.01fF
C11263 VDD3V3 AMUX4_3V_0|SEL[1] 2.19fF
C11264 VDD3V3 BU_3VX2_51|Q 0.16fF
C11265 LS_3VX2_21|Q BU_3VX2_43|Q 0.40fF
C11266 raven_padframe_0|CORNERESDF_3|GNDR raven_padframe_0|CORNERESDF_3|GNDO 0.81fF
C11267 BU_3VX2_23|A BU_3VX2_8|A 0.01fF
C11268 BU_3VX2_10|A BU_3VX2_37|A 0.81fF
C11269 BU_3VX2_0|A BU_3VX2_16|A 0.16fF
C11270 raven_padframe_0|FILLER20F_6|VDDR raven_padframe_0|FILLER20F_6|VDDO 0.06fF
C11271 BU_3VX2_0|A BU_3VX2_29|A 0.01fF
C11272 BU_3VX2_17|A BU_3VX2_31|A 0.01fF
C11273 LS_3VX2_6|Q LS_3VX2_24|Q 0.01fF
C11274 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<14> 33.74fF
C11275 BU_3VX2_63|Q BU_3VX2_0|Q 104.15fF
C11276 raven_padframe_0|CORNERESDF_1|VDDO raven_padframe_0|CORNERESDF_1|GNDO 2.28fF
C11277 raven_soc_0|flash_io2_di BU_3VX2_33|Q 0.01fF
C11278 AMUX4_3V_3|SEL[1] vdd 4.08fF
C11279 AMUX4_3V_1|SEL[0] BU_3VX2_53|Q 63.26fF
C11280 LS_3VX2_27|A BU_3VX2_42|Q 56.66fF
C11281 raven_soc_0|ram_wdata<26> apllc03_1v8_0|CLK 0.01fF
C11282 BU_3VX2_35|A BU_3VX2_5|A 1.21fF
C11283 BU_3VX2_37|A BU_3VX2_0|A 0.01fF
C11284 LS_3VX2_12|A LS_3VX2_6|A 32.27fF
C11285 LS_3VX2_8|Q LS_3VX2_24|Q 0.01fF
C11286 raven_soc_0|gpio_pulldown<0> BU_3VX2_63|Q 0.01fF
C11287 raven_soc_0|gpio_in<0> raven_soc_0|gpio_outenb<10> 0.01fF
C11288 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<14> 0.01fF
C11289 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pulldown<15> 0.01fF
C11290 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_out<13> 19.71fF
C11291 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_out<11> 144.46fF
C11292 raven_soc_0|gpio_out<5> raven_soc_0|gpio_out<7> 1.27fF
C11293 BU_3VX2_20|A raven_soc_0|ext_clk 0.01fF
C11294 LS_3VX2_7|Q VDD3V3 0.16fF
C11295 BU_3VX2_66|A VDD3V3 0.02fF
C11296 BU_3VX2_0|Q raven_soc_0|ram_wdata<16> 0.02fF
C11297 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<31> 5.49fF
C11298 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<1> 1.26fF
C11299 raven_soc_0|flash_io3_di raven_soc_0|flash_io0_di 93.80fF
C11300 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<15> 6.09fF
C11301 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<13> 0.03fF
C11302 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<16> 42.98fF
C11303 raven_soc_0|flash_io1_di raven_soc_0|flash_io1_oeb 17.89fF
C11304 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<31> 3.69fF
C11305 raven_soc_0|ram_wdata<23> raven_soc_0|ram_addr<0> 0.01fF
C11306 raven_soc_0|ram_rdata<30> raven_soc_0|ram_rdata<17> 5.19fF
C11307 LS_3VX2_16|A BU_3VX2_59|Q 22.23fF
C11308 BU_3VX2_41|A BU_3VX2_44|Q 0.02fF
C11309 raven_padframe_0|ICFC_0|GNDR raven_padframe_0|ICFC_0|VDDO 0.09fF
C11310 raven_padframe_0|FILLER20F_2|GNDR raven_padframe_0|FILLER20F_2|GNDO 0.81fF
C11311 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<11> 0.56fF
C11312 BU_3VX2_24|A vdd 0.06fF
C11313 BU_3VX2_38|A raven_soc_0|flash_clk 0.01fF
C11314 BU_3VX2_19|A raven_soc_0|flash_io2_oeb 0.01fF
C11315 VDD BU_3VX2_28|Q 0.05fF
C11316 raven_padframe_0|VDDPADFC_0|VDDR raven_padframe_0|VDDPADFC_0|VDDO 0.06fF
C11317 LS_3VX2_14|A BU_3VX2_62|Q 0.02fF
C11318 BU_3VX2_31|A raven_soc_0|gpio_pulldown<7> 0.01fF
C11319 raven_soc_0|gpio_in<4> VDD3V3 0.24fF
C11320 VDD raven_padframe_0|CORNERESDF_0|GNDO 0.07fF
C11321 AMUX2_3V_0|SEL BU_3VX2_57|Q 0.01fF
C11322 raven_soc_0|gpio_pullup<9> BU_3VX2_26|Q 0.01fF
C11323 BU_3VX2_9|A BU_3VX2_38|A 0.76fF
C11324 BU_3VX2_6|A BU_3VX2_19|A 0.84fF
C11325 BU_3VX2_10|A LS_3VX2_3|Q 3.37fF
C11326 LS_3VX2_14|A LS_3VX2_5|A 11.13fF
C11327 BU_3VX2_31|A BU_3VX2_12|A 0.01fF
C11328 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<6> 1.19fF
C11329 raven_soc_0|gpio_out<4> raven_soc_0|gpio_pullup<4> 0.51fF
C11330 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<10> 1.33fF
C11331 LS_3VX2_3|A raven_soc_0|gpio_pulldown<4> 0.01fF
C11332 BU_3VX2_25|A raven_soc_0|flash_io3_do 0.01fF
C11333 BU_3VX2_63|Q raven_soc_0|flash_io3_di 0.01fF
C11334 IN_3VX2_1|A LS_3VX2_21|A 0.01fF
C11335 BU_3VX2_14|A raven_soc_0|flash_io2_di 0.01fF
C11336 raven_soc_0|ext_clk raven_soc_0|gpio_in<13> 0.18fF
C11337 BU_3VX2_40|Q raven_soc_0|gpio_in<8> 0.01fF
C11338 raven_soc_0|gpio_in<7> VDD3V3 0.07fF
C11339 raven_soc_0|gpio_pullup<5> raven_soc_0|gpio_in<9> 0.02fF
C11340 BU_3VX2_55|A BU_3VX2_56|A 10.09fF
C11341 BU_3VX2_52|A BU_3VX2_59|A 0.50fF
C11342 BU_3VX2_54|A BU_3VX2_57|A 1.72fF
C11343 BU_3VX2_53|A BU_3VX2_58|A 0.84fF
C11344 VDD3V3 BU_3VX2_61|A 0.10fF
C11345 LS_3VX2_8|Q LS_3VX2_6|Q 1.80fF
C11346 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<0> 21.25fF
C11347 BU_3VX2_0|A LS_3VX2_3|Q 0.01fF
C11348 BU_3VX2_8|A IN_3VX2_1|A 0.01fF
C11349 IN_3VX2_1|A raven_soc_0|gpio_pulldown<1> 0.01fF
C11350 LOGIC0_3V_4|Q raven_soc_0|gpio_pulldown<12> 0.01fF
C11351 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pullup<12> 0.02fF
C11352 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_in<3> 1.78fF
C11353 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<5> 0.02fF
C11354 raven_spi_0|sdo_enb raven_soc_0|gpio_pullup<15> 1.01fF
C11355 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<10> 0.01fF
C11356 raven_soc_0|gpio_out<2> BU_3VX2_0|Q 0.01fF
C11357 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<8> 0.01fF
C11358 raven_soc_0|ram_wdata<4> raven_soc_0|ram_rdata<19> 0.04fF
C11359 raven_soc_0|gpio_pullup<13> BU_3VX2_40|Q 0.02fF
C11360 raven_soc_0|gpio_pulldown<6> raven_soc_0|gpio_in<12> 0.02fF
C11361 raven_soc_0|flash_io0_di raven_soc_0|irq_pin 0.01fF
C11362 raven_soc_0|irq_pin BU_3VX2_46|Q 13.12fF
C11363 BU_3VX2_66|Q BU_3VX2_24|Q 1.35fF
C11364 BU_3VX2_19|Q BU_3VX2_27|Q 9.93fF
C11365 BU_3VX2_38|Q BU_3VX2_28|Q 0.14fF
C11366 BU_3VX2_2|Q BU_3VX2_23|Q 2.18fF
C11367 BU_3VX2_21|Q BU_3VX2_25|Q 9.48fF
C11368 BU_3VX2_15|Q BU_3VX2_29|Q 0.01fF
C11369 BU_3VX2_67|Q BU_3VX2_28|Q 0.06fF
C11370 BU_3VX2_18|Q BU_3VX2_27|Q 11.00fF
C11371 BU_3VX2_8|Q BU_3VX2_25|Q 0.81fF
C11372 BU_3VX2_9|Q BU_3VX2_29|Q 1.39fF
C11373 BU_3VX2_20|Q BU_3VX2_24|Q 9.46fF
C11374 LS_3VX2_17|A BU_3VX2_53|Q 7.85fF
C11375 BU_3VX2_10|Q BU_3VX2_23|Q 2.85fF
C11376 BU_3VX2_61|Q BU_3VX2_57|Q 34.96fF
C11377 LS_3VX2_15|A BU_3VX2_55|Q 13.90fF
C11378 AMUX4_3V_4|AIN2 BU_3VX2_52|Q 0.01fF
C11379 BU_3VX2_22|Q apllc03_1v8_0|CLK 0.01fF
C11380 BU_3VX2_17|Q BU_3VX2_26|Q 3.87fF
C11381 BU_3VX2_62|Q BU_3VX2_56|Q 19.44fF
C11382 BU_3VX2_22|A BU_3VX2_17|A 3.82fF
C11383 LS_3VX2_8|A LS_3VX2_13|A 150.32fF
C11384 raven_soc_0|gpio_pulldown<0> raven_soc_0|gpio_out<2> 8.79fF
C11385 raven_soc_0|gpio_in<4> raven_soc_0|gpio_outenb<6> 0.87fF
C11386 LS_3VX2_5|A BU_3VX2_56|Q 18.80fF
C11387 BU_3VX2_0|Q BU_3VX2_68|Q 0.01fF
C11388 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_out<8> 22.33fF
C11389 AMUX4_3V_3|SEL[1] BU_3VX2_70|Q 2.26fF
C11390 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<18> 19.81fF
C11391 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<5> 0.04fF
C11392 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<21> 0.32fF
C11393 raven_soc_0|ram_rdata<19> vdd 0.47fF
C11394 raven_soc_0|flash_clk BU_3VX2_23|Q 0.01fF
C11395 raven_soc_0|flash_io1_oeb BU_3VX2_28|Q 11.09fF
C11396 BU_3VX2_41|A vdd 0.06fF
C11397 raven_padframe_0|FILLER50F_0|VDDO raven_padframe_0|FILLER50F_0|GNDO 2.28fF
C11398 raven_padframe_0|aregc01_3v3_1|VDDO raven_padframe_0|aregc01_3v3_1|GNDO 1.69fF
C11399 raven_padframe_0|axtoc02_3v3_0|m4_55000_29333# raven_padframe_0|axtoc02_3v3_0|GNDO 0.25fF
C11400 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<6> 1.04fF
C11401 BU_3VX2_10|A raven_soc_0|flash_io1_oeb 0.01fF
C11402 AMUX4_3V_1|AIN1 BU_3VX2_62|Q 0.14fF
C11403 BU_3VX2_63|A raven_soc_0|flash_io0_di 0.01fF
C11404 BU_3VX2_16|A vdd 0.06fF
C11405 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<15> 0.02fF
C11406 BU_3VX2_29|A vdd 0.06fF
C11407 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_in<12> 14.27fF
C11408 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_in<14> 215.12fF
C11409 raven_soc_0|gpio_outenb<12> raven_soc_0|gpio_in<9> 0.38fF
C11410 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_in<8> 4.37fF
C11411 LS_3VX2_3|A raven_soc_0|flash_io2_di 0.01fF
C11412 adc_low AMUX4_3V_4|AIN2 0.07fF
C11413 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<10> 44.15fF
C11414 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<15> 114.94fF
C11415 raven_soc_0|gpio_outenb<10> raven_soc_0|gpio_in<13> 0.02fF
C11416 raven_soc_0|gpio_out<5> BU_3VX2_40|Q 0.01fF
C11417 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_in<7> 1.88fF
C11418 raven_soc_0|gpio_out<7> VDD3V3 0.07fF
C11419 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<23> 4.84fF
C11420 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<11> 75.19fF
C11421 raven_soc_0|ram_wdata<24> raven_soc_0|ram_rdata<20> 0.02fF
C11422 raven_soc_0|ram_wdata<7> raven_soc_0|ram_rdata<0> 0.01fF
C11423 raven_soc_0|ram_rdata<6> raven_soc_0|ram_rdata<19> 1.97fF
C11424 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<8> 0.01fF
C11425 BU_3VX2_7|A BU_3VX2_18|A 1.03fF
C11426 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<10> 0.01fF
C11427 BU_3VX2_38|A BU_3VX2_28|A 0.01fF
C11428 BU_3VX2_37|A vdd 0.25fF
C11429 BU_3VX2_5|A raven_soc_0|flash_io3_di 0.03fF
C11430 BU_3VX2_0|A raven_soc_0|flash_io1_oeb 3.76fF
C11431 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<3> 19.48fF
C11432 LOGIC0_3V_4|Q comp_inp 1.85fF
C11433 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_pullup<14> 13.72fF
C11434 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<13> 0.07fF
C11435 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<10> 0.09fF
C11436 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_pullup<13> 0.02fF
C11437 raven_soc_0|gpio_outenb<0> BU_3VX2_71|Q 0.01fF
C11438 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_pullup<6> 0.02fF
C11439 raven_soc_0|gpio_out<6> raven_soc_0|gpio_pulldown<7> 1.78fF
C11440 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<5> 0.05fF
C11441 AMUX2_3V_0|SEL LS_3VX2_16|A 0.01fF
C11442 raven_padframe_0|BBCUD4F_6|VDDR raven_padframe_0|BBCUD4F_6|GNDO 0.13fF
C11443 raven_soc_0|gpio_pulldown<15> BU_3VX2_24|Q 0.01fF
C11444 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<12> 0.02fF
C11445 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<15> 3.04fF
C11446 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<8> 0.71fF
C11447 BU_3VX2_16|Q BU_3VX2_68|Q 0.04fF
C11448 BU_3VX2_64|Q BU_3VX2_69|Q 6.53fF
C11449 BU_3VX2_68|Q BU_3VX2_30|Q 0.49fF
C11450 VDD3V3 BU_3VX2_49|Q 0.14fF
C11451 LS_3VX2_20|Q BU_3VX2_42|Q 5.34fF
C11452 BU_3VX2_22|A BU_3VX2_12|A 1.53fF
C11453 BU_3VX2_3|A BU_3VX2_26|A 0.01fF
C11454 BU_3VX2_40|A BU_3VX2_29|A 0.13fF
C11455 BU_3VX2_19|A BU_3VX2_27|A 2.65fF
C11456 BU_3VX2_63|A BU_3VX2_63|Q 0.08fF
C11457 BU_3VX2_15|A BU_3VX2_26|A 1.86fF
C11458 LS_3VX2_8|A raven_soc_0|ser_rx 0.01fF
C11459 raven_soc_0|gpio_pulldown<11> LS_3VX2_3|A 0.01fF
C11460 LS_3VX2_4|A LS_3VX2_13|A 9.16fF
C11461 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_1|PO 0.04fF
C11462 AMUX4_3V_1|SEL[1] BU_3VX2_55|Q 21.87fF
C11463 raven_soc_0|ram_wdata<28> apllc03_1v8_0|CLK 0.01fF
C11464 raven_soc_0|gpio_in<1> raven_soc_0|gpio_in<3> 4.45fF
C11465 BU_3VX2_56|Q BU_3VX2_45|Q 0.16fF
C11466 raven_soc_0|gpio_in<1> raven_soc_0|gpio_out<9> 0.09fF
C11467 BU_3VX2_8|A BU_3VX2_25|A 0.01fF
C11468 BU_3VX2_37|A BU_3VX2_40|A 5.43fF
C11469 BU_3VX2_21|A BU_3VX2_17|A 4.96fF
C11470 BU_3VX2_3|A BU_3VX2_11|A 1.24fF
C11471 raven_soc_0|gpio_out<0> IN_3VX2_1|A 0.01fF
C11472 BU_3VX2_15|A BU_3VX2_11|A 4.87fF
C11473 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pullup<10> 0.01fF
C11474 IN_3VX2_1|A raven_soc_0|gpio_out<12> 0.01fF
C11475 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_out<11> 22.44fF
C11476 raven_soc_0|gpio_outenb<14> raven_soc_0|gpio_outenb<15> 31.93fF
C11477 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_out<9> 0.63fF
C11478 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_out<7> 3.87fF
C11479 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<5> 0.45fF
C11480 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_out<13> 0.01fF
C11481 raven_soc_0|gpio_outenb<7> raven_soc_0|gpio_out<5> 0.02fF
C11482 LS_3VX2_4|Q VDD3V3 0.16fF
C11483 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pullup<5> 0.19fF
C11484 LS_3VX2_7|A BU_3VX2_55|Q 6.86fF
C11485 raven_soc_0|gpio_outenb<1> raven_soc_0|ext_clk 0.15fF
C11486 raven_soc_0|ram_addr<7> raven_soc_0|ram_addr<3> 15.63fF
C11487 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<31> 26.29fF
C11488 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<6> 0.35fF
C11489 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<23> 0.01fF
C11490 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<20> 0.01fF
C11491 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<30> 4.91fF
C11492 raven_soc_0|ram_wdata<24> raven_soc_0|ram_wdata<17> 10.97fF
C11493 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<13> 0.39fF
C11494 raven_soc_0|ram_rdata<7> raven_soc_0|ram_rdata<17> 4.77fF
C11495 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<29> 16.07fF
C11496 BU_3VX2_12|Q BU_3VX2_36|Q 5.90fF
C11497 BU_3VX2_2|Q BU_3VX2_4|Q 27.23fF
C11498 BU_3VX2_4|Q BU_3VX2_10|Q 12.02fF
C11499 raven_soc_0|flash_io1_do raven_soc_0|flash_io2_di 59.53fF
C11500 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<27> 2.67fF
C11501 BU_3VX2_11|Q BU_3VX2_17|Q 6.19fF
C11502 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<1> 0.18fF
C11503 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<31> 0.02fF
C11504 raven_soc_0|ram_rdata<10> raven_soc_0|ram_rdata<2> 2.68fF
C11505 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<19> 0.01fF
C11506 raven_soc_0|ram_addr<2> raven_soc_0|ram_wdata<21> 0.01fF
C11507 raven_soc_0|ram_addr<4> raven_soc_0|ram_wdata<25> 0.01fF
C11508 LOGIC0_3V_0|Q LOGIC0_3V_4|Q 0.01fF
C11509 LS_3VX2_16|A BU_3VX2_61|Q 36.13fF
C11510 AMUX4_3V_4|AIN2 BU_3VX2_58|Q 0.01fF
C11511 raven_spi_0|SDO raven_soc_0|flash_io0_di 2.27fF
C11512 BU_3VX2_2|A raven_soc_0|flash_io3_oeb 0.01fF
C11513 raven_soc_0|gpio_in<1> raven_padframe_0|BBCUD4F_0|PO 0.04fF
C11514 BU_3VX2_4|A raven_soc_0|flash_io3_do 0.01fF
C11515 LS_3VX2_11|A BU_3VX2_54|Q 8.41fF
C11516 LS_3VX2_3|Q vdd 0.24fF
C11517 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pulldown<7> 0.28fF
C11518 AMUX2_3V_0|AOUT AMUX4_3V_4|AIN2 0.32fF
C11519 raven_soc_0|gpio_pulldown<13> BU_3VX2_28|Q 0.01fF
C11520 BU_3VX2_0|Q BU_3VX2_24|Q 0.02fF
C11521 raven_soc_0|gpio_pulldown<9> BU_3VX2_26|Q 0.01fF
C11522 BU_3VX2_71|Q raven_soc_0|flash_io0_do 0.08fF
C11523 BU_3VX2_68|A BU_3VX2_1|A 0.54fF
C11524 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pulldown<12> 31.83fF
C11525 LS_3VX2_4|A raven_soc_0|ser_rx 0.01fF
C11526 AMUX4_3V_4|AOUT AMUX4_3V_4|AIN3 10.70fF
C11527 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<15> 0.91fF
C11528 LOGIC0_3V_4|Q vdd 2.11fF
C11529 IN_3VX2_1|A LS_3VX2_27|A 0.01fF
C11530 raven_soc_0|gpio_pulldown<0> BU_3VX2_24|Q 0.01fF
C11531 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<15> 67.87fF
C11532 raven_soc_0|gpio_pullup<1> BU_3VX2_28|Q 0.01fF
C11533 raven_soc_0|gpio_outenb<2> BU_3VX2_29|Q 0.01fF
C11534 BU_3VX2_40|Q VDD3V3 0.06fF
C11535 LS_3VX2_21|Q LS_3VX2_27|Q 13.70fF
C11536 LS_3VX2_20|Q BU_3VX2_42|A 2.05fF
C11537 VDD raven_padframe_0|FILLER50F_2|VDDR 0.71fF
C11538 LS_3VX2_9|A LS_3VX2_10|A 54.55fF
C11539 BU_3VX2_7|A BU_3VX2_71|A 0.02fF
C11540 BU_3VX2_63|A BU_3VX2_5|A 0.01fF
C11541 LS_3VX2_3|Q BU_3VX2_40|A 0.01fF
C11542 BU_3VX2_21|A BU_3VX2_12|A 1.73fF
C11543 raven_padframe_0|BBCUD4F_3|GNDR raven_padframe_0|BBCUD4F_3|VDDO 0.09fF
C11544 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pullup<3> 1.81fF
C11545 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<0> 0.29fF
C11546 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_outenb<10> 0.01fF
C11547 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_pulldown<12> 0.01fF
C11548 markings_0|product_name_0|_alphabet_V_0|m2_0_560# markings_0|product_name_0|_alphabet_A_0|m2_0_0# 0.96fF
C11549 raven_padframe_0|BBCUD4F_14|VDDR raven_padframe_0|BBCUD4F_14|GNDR 0.68fF
C11550 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<5> 0.01fF
C11551 raven_soc_0|gpio_pulldown<14> BU_3VX2_71|Q 0.01fF
C11552 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_6|PO 0.04fF
C11553 raven_soc_0|gpio_pulldown<3> raven_soc_0|ext_clk 0.01fF
C11554 LS_3VX2_22|A AMUX4_3V_4|AIN2 1.73fF
C11555 BU_3VX2_38|Q vdd 1.12fF
C11556 BU_3VX2_19|Q BU_3VX2_25|Q 17.75fF
C11557 BU_3VX2_16|Q BU_3VX2_24|Q 4.43fF
C11558 BU_3VX2_18|Q BU_3VX2_25|Q 13.41fF
C11559 BU_3VX2_64|Q BU_3VX2_29|Q 0.01fF
C11560 BU_3VX2_67|Q vdd 0.91fF
C11561 VDD3V3 raven_padframe_0|VDDORPADF_4|GNDO 2.41fF
C11562 BU_3VX2_65|Q BU_3VX2_28|Q 0.26fF
C11563 BU_3VX2_30|Q BU_3VX2_24|Q 5.37fF
C11564 LS_3VX2_15|A BU_3VX2_57|Q 20.18fF
C11565 BU_3VX2_31|Q apllc03_1v8_0|CLK 3.75fF
C11566 raven_soc_0|gpio_in<9> raven_padframe_0|BBCUD4F_9|PO 0.04fF
C11567 raven_spi_0|CSB raven_spi_0|sdo_enb 33.27fF
C11568 raven_padframe_0|FILLER50F_2|VDDR LOGIC0_3V_4|Q 0.01fF
C11569 LOGIC0_3V_4|Q raven_soc_0|gpio_in<2> 0.54fF
C11570 LS_3VX2_14|Q LS_3VX2_24|Q 0.45fF
C11571 raven_soc_0|gpio_in<4> raven_soc_0|gpio_pullup<8> 0.01fF
C11572 raven_soc_0|gpio_pulldown<7> raven_soc_0|gpio_pulldown<6> 16.03fF
C11573 raven_soc_0|ram_rdata<1> raven_soc_0|ram_rdata<17> 1.12fF
C11574 raven_soc_0|ram_wdata<27> raven_soc_0|ram_rdata<15> 0.54fF
C11575 raven_soc_0|ram_wdata<31> raven_soc_0|ram_addr<0> 0.02fF
C11576 raven_soc_0|flash_io1_oeb vdd 2.29fF
C11577 BU_3VX2_58|A BU_3VX2_58|Q 0.10fF
C11578 raven_soc_0|flash_io0_di BU_3VX2_26|Q 0.01fF
C11579 raven_soc_0|flash_io2_oeb BU_3VX2_27|Q 0.01fF
C11580 raven_soc_0|flash_io3_oeb apllc03_1v8_0|CLK 0.01fF
C11581 raven_soc_0|flash_io3_di BU_3VX2_24|Q 0.01fF
C11582 adc0_data<5> BU_3VX2_51|Q 26.95fF
C11583 AMUX4_3V_0|SEL[1] adc0_data<5> 20.00fF
C11584 raven_padframe_0|FILLER01F_1|VDDR raven_padframe_0|FILLER01F_1|VDDO 0.06fF
C11585 raven_padframe_0|BBC4F_3|GNDR raven_padframe_0|BBC4F_3|GNDO 0.81fF
C11586 raven_padframe_0|VDDORPADF_4|GNDR raven_padframe_0|VDDORPADF_4|GNDO 0.81fF
C11587 raven_padframe_0|axtoc02_3v3_0|m4_55000_28769# raven_padframe_0|axtoc02_3v3_0|m4_55000_22024# 0.06fF
C11588 raven_soc_0|gpio_out<3> raven_soc_0|gpio_out<13> 0.01fF
C11589 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_out<11> 4.13fF
C11590 raven_soc_0|gpio_in<1> raven_soc_0|ext_clk 0.01fF
C11591 BU_3VX2_3|A VDD3V3 0.20fF
C11592 BU_3VX2_15|A VDD3V3 0.48fF
C11593 raven_soc_0|gpio_outenb<6> BU_3VX2_40|Q 1.69fF
C11594 BU_3VX2_0|Q raven_soc_0|gpio_out<15> 0.07fF
C11595 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_in<14> 18.82fF
C11596 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_in<13> 5.88fF
C11597 raven_soc_0|gpio_pullup<12> raven_soc_0|gpio_in<9> 0.01fF
C11598 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_in<12> 34.05fF
C11599 raven_soc_0|gpio_outenb<7> VDD3V3 0.07fF
C11600 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_in<6> 2.15fF
C11601 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_in<8> 6.32fF
C11602 raven_soc_0|gpio_outenb<5> raven_soc_0|ext_clk 0.01fF
C11603 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_in<7> 4.23fF
C11604 raven_soc_0|ser_rx comp_inp 33.65fF
C11605 raven_soc_0|ram_rdata<4> raven_soc_0|ram_rdata<0> 4.69fF
C11606 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<20> 5.28fF
C11607 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<23> 15.87fF
C11608 raven_soc_0|ram_rdata<24> raven_soc_0|ram_rdata<19> 22.94fF
C11609 raven_soc_0|ram_addr<3> raven_soc_0|ram_rdata<11> 2.85fF
C11610 raven_spi_0|CSB raven_soc_0|gpio_in<15> 1.84fF
C11611 BU_3VX2_38|A LS_3VX2_3|A 0.52fF
C11612 BU_3VX2_40|A raven_soc_0|flash_io1_oeb 0.01fF
C11613 BU_3VX2_31|A raven_soc_0|flash_clk 65.27fF
C11614 LOGIC0_3V_4|Q raven_soc_0|gpio_in<11> 0.08fF
C11615 BU_3VX2_13|A raven_soc_0|flash_io3_di 0.01fF
C11616 BU_3VX2_0|Q raven_soc_0|gpio_in<5> 0.01fF
C11617 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<3> 0.26fF
C11618 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_pullup<13> 0.91fF
C11619 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<14> 0.57fF
C11620 raven_soc_0|ram_wenb raven_soc_0|ram_rdata<26> 0.07fF
C11621 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_pullup<6> 0.02fF
C11622 raven_soc_0|gpio_outenb<11> raven_soc_0|gpio_pulldown<7> 0.02fF
C11623 raven_soc_0|gpio_pulldown<10> BU_3VX2_71|Q 0.01fF
C11624 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<14> 0.02fF
C11625 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<10> 3.32fF
C11626 BU_3VX2_33|A raven_soc_0|flash_io0_oeb 0.01fF
C11627 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<13> 0.02fF
C11628 BU_3VX2_0|Q LS_3VX2_23|A 0.37fF
C11629 raven_soc_0|gpio_outenb<4> apllc03_1v8_0|CLK 0.01fF
C11630 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<14> 2.25fF
C11631 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<15> 2.60fF
C11632 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<13> 0.01fF
C11633 LS_3VX2_13|A vdd 2.38fF
C11634 BU_3VX2_63|Q BU_3VX2_26|Q 2.10fF
C11635 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<9> 10.24fF
C11636 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<1> 7.20fF
C11637 raven_soc_0|ram_wdata<9> raven_soc_0|ram_wdata<0> 2.12fF
C11638 raven_soc_0|ram_wdata<0> raven_soc_0|ram_wdata<1> 40.12fF
C11639 BU_3VX2_8|A BU_3VX2_4|A 3.22fF
C11640 LS_3VX2_11|A LS_3VX2_14|A 18.69fF
C11641 BU_3VX2_9|A BU_3VX2_31|A 0.01fF
C11642 LS_3VX2_6|Q LS_3VX2_14|Q 0.58fF
C11643 raven_padframe_0|VDDPADF_0|GNDR raven_padframe_0|VDDPADF_0|GNDO 0.81fF
C11644 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<9> 0.01fF
C11645 raven_padframe_0|BT4F_0|VDDR raven_padframe_0|BT4F_0|VDDO 0.06fF
C11646 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_8|PO 0.04fF
C11647 AMUX4_3V_1|SEL[1] BU_3VX2_57|Q 15.87fF
C11648 raven_soc_0|ram_wdata<15> vdd 0.76fF
C11649 raven_soc_0|gpio_in<1> raven_soc_0|gpio_outenb<10> 0.01fF
C11650 LS_3VX2_8|Q LS_3VX2_14|Q 0.31fF
C11651 raven_spi_0|SDI LOGIC0_3V_3|Q 2.39fF
C11652 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pullup<3> 0.01fF
C11653 IN_3VX2_1|A raven_soc_0|gpio_outenb<12> 0.01fF
C11654 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<14> 0.01fF
C11655 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<4> 0.01fF
C11656 raven_soc_0|gpio_pullup<15> raven_soc_0|gpio_outenb<15> 69.44fF
C11657 raven_soc_0|gpio_outenb<6> raven_soc_0|gpio_outenb<7> 11.02fF
C11658 raven_soc_0|gpio_outenb<5> raven_soc_0|gpio_outenb<10> 0.83fF
C11659 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pullup<7> 0.01fF
C11660 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_out<5> 0.01fF
C11661 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_out<9> 6.31fF
C11662 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_out<7> 3.13fF
C11663 LS_3VX2_7|A BU_3VX2_57|Q 0.01fF
C11664 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<26> 2.39fF
C11665 BU_3VX2_2|Q BU_3VX2_3|Q 78.33fF
C11666 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<4> 5.44fF
C11667 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<15> 0.07fF
C11668 raven_soc_0|ram_wdata<16> raven_soc_0|ram_rdata<10> 0.12fF
C11669 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<30> 37.81fF
C11670 BU_3VX2_15|Q BU_3VX2_32|Q 0.15fF
C11671 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<4> 0.32fF
C11672 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<9> 3.44fF
C11673 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<24> 14.11fF
C11674 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<23> 0.12fF
C11675 raven_soc_0|ram_rdata<10> raven_soc_0|ram_wdata<2> 0.09fF
C11676 BU_3VX2_38|Q BU_3VX2_70|Q 0.85fF
C11677 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<19> 0.02fF
C11678 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<21> 0.02fF
C11679 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<25> 2.41fF
C11680 raven_soc_0|ram_rdata<7> raven_soc_0|ram_wdata<22> 0.02fF
C11681 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<17> 0.01fF
C11682 raven_soc_0|ram_rdata<3> raven_soc_0|ram_addr<2> 0.04fF
C11683 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<21> 0.01fF
C11684 raven_soc_0|flash_io3_do raven_soc_0|flash_io0_oeb 19.12fF
C11685 AMUX4_3V_3|SEL[1] LS_3VX2_2|A 1.53fF
C11686 BU_3VX2_36|Q BU_3VX2_5|Q 2.14fF
C11687 BU_3VX2_32|Q BU_3VX2_9|Q 8.85fF
C11688 BU_3VX2_70|Q BU_3VX2_67|Q 6.75fF
C11689 BU_3VX2_3|Q BU_3VX2_10|Q 6.59fF
C11690 BU_3VX2_37|Q BU_3VX2_8|Q 5.26fF
C11691 raven_soc_0|flash_io0_oeb AMUX4_3V_4|AIN3 2.34fF
C11692 AMUX4_3V_4|AIN2 BU_3VX2_60|Q 0.01fF
C11693 LS_3VX2_16|A LS_3VX2_15|A 60.57fF
C11694 BU_3VX2_25|Q BU_3VX2_27|Q 114.03fF
C11695 apllc03_1v8_0|B_VCO BU_3VX2_29|Q 0.35fF
C11696 BU_3VX2_23|Q apllc03_1v8_0|B_CP 0.66fF
C11697 raven_padframe_0|BBCUD4F_15|GNDR raven_padframe_0|BBCUD4F_15|GNDO 0.81fF
C11698 BU_3VX2_6|A raven_soc_0|flash_io2_oeb 0.01fF
C11699 AMUX4_3V_1|AIN1 AMUX4_3V_4|AIN3 2.69fF
C11700 BU_3VX2_38|A raven_soc_0|flash_io1_do 0.01fF
C11701 IN_3VX2_1|Q BU_3VX2_55|Q 0.01fF
C11702 LS_3VX2_11|A BU_3VX2_56|Q 11.17fF
C11703 VDD raven_padframe_0|FILLER20F_4|VDDR 0.71fF
C11704 raven_soc_0|gpio_pulldown<13> vdd 0.31fF
C11705 raven_soc_0|ser_rx vdd 5.38fF
C11706 LS_3VX2_3|A BU_3VX2_23|Q 0.01fF
C11707 raven_padframe_0|BBCUD4F_5|VDDR raven_padframe_0|BBCUD4F_5|GNDO 0.13fF
C11708 BU_3VX2_71|Q raven_soc_0|flash_io1_di 0.09fF
C11709 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<15> 0.36fF
C11710 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<16> 18.61fF
C11711 raven_soc_0|gpio_out<1> raven_soc_0|gpio_outenb<2> 11.59fF
C11712 raven_soc_0|gpio_out<4> LS_3VX2_3|A 0.01fF
C11713 LS_3VX2_9|A raven_soc_0|ser_tx 0.01fF
C11714 LS_3VX2_14|A LS_3VX2_21|A 9.65fF
C11715 LS_3VX2_8|A AMUX4_3V_1|SEL[0] 12.89fF
C11716 raven_soc_0|gpio_out<3> raven_soc_0|gpio_in<14> 0.02fF
C11717 VDD raven_padframe_0|APR00DF_1|GNDR 0.16fF
C11718 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<10> 12.37fF
C11719 BU_3VX2_0|Q raven_soc_0|ram_wdata<20> 0.02fF
C11720 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_in<6> 0.01fF
C11721 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_in<12> 0.02fF
C11722 BU_3VX2_27|A BU_3VX2_27|Q 0.08fF
C11723 raven_soc_0|gpio_pullup<1> vdd 0.18fF
C11724 raven_soc_0|gpio_out<2> BU_3VX2_26|Q 0.99fF
C11725 BU_3VX2_24|A BU_3VX2_7|A 0.01fF
C11726 VDD raven_padframe_0|APR00DF_1|VDDR 0.71fF
C11727 LS_3VX2_9|A LS_3VX2_24|A 7.31fF
C11728 BU_3VX2_63|A BU_3VX2_13|A 0.01fF
C11729 BU_3VX2_31|A BU_3VX2_28|A 19.44fF
C11730 raven_soc_0|gpio_pulldown<1> raven_soc_0|gpio_pulldown<5> 1.50fF
C11731 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<10> 0.03fF
C11732 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pulldown<13> 0.01fF
C11733 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pullup<10> 0.71fF
C11734 BU_3VX2_22|A raven_soc_0|flash_clk 1.92fF
C11735 raven_soc_0|gpio_pulldown<2> raven_soc_0|gpio_pullup<4> 6.95fF
C11736 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_outenb<8> 0.66fF
C11737 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<14> 241.50fF
C11738 raven_soc_0|gpio_in<0> raven_soc_0|flash_io2_di 0.26fF
C11739 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pullup<6> 0.01fF
C11740 BU_3VX2_63|Q raven_soc_0|gpio_outenb<13> 0.01fF
C11741 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<10> 0.01fF
C11742 raven_soc_0|flash_csb raven_soc_0|flash_io2_di 13.52fF
C11743 BU_3VX2_65|Q vdd 1.49fF
C11744 BU_3VX2_68|Q BU_3VX2_26|Q 0.01fF
C11745 BU_3VX2_22|A BU_3VX2_9|A 1.58fF
C11746 LS_3VX2_7|Q LS_3VX2_24|Q 0.01fF
C11747 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<1> 21.53fF
C11748 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<0> 10.56fF
C11749 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<31> 0.01fF
C11750 raven_soc_0|ram_addr<6> raven_soc_0|ram_rdata<17> 0.01fF
C11751 raven_soc_0|ram_wdata<29> raven_soc_0|ram_wdata<31> 69.10fF
C11752 raven_soc_0|ram_wdata<22> raven_soc_0|ram_rdata<1> 1.51fF
C11753 raven_soc_0|ram_wdata<25> raven_soc_0|ram_rdata<13> 0.02fF
C11754 raven_soc_0|ram_wdata<26> raven_soc_0|ram_rdata<15> 0.44fF
C11755 raven_soc_0|ram_wdata<19> raven_soc_0|ram_addr<0> 0.01fF
C11756 raven_soc_0|ram_wdata<17> raven_soc_0|ram_rdata<16> 0.01fF
C11757 AMUX4_3V_1|SEL[1] LS_3VX2_16|A 0.12fF
C11758 BU_3VX2_56|Q LS_3VX2_21|A 0.03fF
C11759 BU_3VX2_47|A BU_3VX2_42|A 0.18fF
C11760 BU_3VX2_41|A LS_3VX2_21|Q 0.21fF
C11761 BU_3VX2_46|A BU_3VX2_43|A 0.83fF
C11762 BU_3VX2_45|A BU_3VX2_44|A 5.87fF
C11763 raven_soc_0|flash_io1_do BU_3VX2_23|Q 0.01fF
C11764 raven_soc_0|flash_io3_do BU_3VX2_29|Q 0.01fF
C11765 raven_soc_0|flash_io2_oeb BU_3VX2_25|Q 0.01fF
C11766 LS_3VX2_16|Q BU_3VX2_61|Q 0.40fF
C11767 BU_3VX2_58|A BU_3VX2_60|Q 0.03fF
C11768 AMUX4_3V_0|SEL[0] BU_3VX2_46|Q 18.90fF
C11769 adc0_data<5> BU_3VX2_49|Q 47.19fF
C11770 BU_3VX2_44|Q BU_3VX2_72|Q 1.02fF
C11771 raven_soc_0|gpio_pullup<2> LOGIC0_3V_4|Q 0.06fF
C11772 raven_soc_0|gpio_out<3> raven_soc_0|gpio_outenb<15> 0.49fF
C11773 raven_soc_0|gpio_in<3> raven_soc_0|gpio_pulldown<15> 0.01fF
C11774 raven_soc_0|gpio_in<0> raven_soc_0|gpio_pulldown<11> 0.01fF
C11775 raven_padframe_0|axtoc02_3v3_0|m4_55000_30133# raven_padframe_0|axtoc02_3v3_0|m4_55000_29057# 0.02fF
C11776 raven_padframe_0|axtoc02_3v3_0|m4_0_30653# raven_padframe_0|axtoc02_3v3_0|VDDR 0.15fF
C11777 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_out<9> 0.01fF
C11778 markings_0|date_0|_alphabet_0_0|m2_0_208# markings_0|date_0|_alphabet_2_0|m2_0_0# 0.69fF
C11779 raven_spi_0|SDI VDD3V3 1.73fF
C11780 raven_padframe_0|POWERCUTVDD3FC_0|VDDR raven_padframe_0|POWERCUTVDD3FC_0|GNDO 0.13fF
C11781 LS_3VX2_7|A LS_3VX2_16|A 0.01fF
C11782 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_in<11> 7.81fF
C11783 LS_3VX2_4|A AMUX4_3V_1|SEL[0] 55.59fF
C11784 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_in<9> 0.22fF
C11785 raven_soc_0|gpio_pullup<8> BU_3VX2_40|Q 0.02fF
C11786 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<5> 1.00fF
C11787 adc_high BU_3VX2_53|Q 0.30fF
C11788 raven_soc_0|gpio_pullup<7> raven_soc_0|ext_clk 0.01fF
C11789 raven_soc_0|gpio_pullup<9> VDD3V3 0.07fF
C11790 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_in<8> 7.45fF
C11791 BU_3VX2_0|Q raven_soc_0|gpio_in<6> 0.01fF
C11792 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<11> 0.01fF
C11793 raven_soc_0|ram_rdata<22> raven_soc_0|ram_rdata<20> 48.68fF
C11794 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<28> 11.63fF
C11795 BU_3VX2_71|Q BU_3VX2_28|Q 2.72fF
C11796 raven_soc_0|gpio_outenb<8> apllc03_1v8_0|CLK 0.01fF
C11797 raven_soc_0|gpio_out<14> BU_3VX2_29|Q 0.01fF
C11798 BU_3VX2_36|Q BU_3VX2_28|Q 14.23fF
C11799 BU_3VX2_8|A raven_soc_0|flash_io0_oeb 0.01fF
C11800 BU_3VX2_20|A raven_soc_0|flash_io2_di 0.01fF
C11801 LS_3VX2_8|A LS_3VX2_17|A 0.01fF
C11802 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pulldown<6> 0.39fF
C11803 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<9> 7.13fF
C11804 BU_3VX2_0|Q raven_soc_0|gpio_out<10> 0.48fF
C11805 BU_3VX2_33|A raven_soc_0|flash_io2_do 0.20fF
C11806 raven_soc_0|gpio_pulldown<12> BU_3VX2_71|Q 0.01fF
C11807 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<9> 0.01fF
C11808 raven_soc_0|gpio_pullup<11> raven_soc_0|gpio_pulldown<7> 0.02fF
C11809 raven_soc_0|ram_wdata<3> raven_soc_0|ram_wdata<11> 3.22fF
C11810 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_pullup<14> 0.02fF
C11811 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<13> 0.02fF
C11812 BU_3VX2_27|A raven_soc_0|flash_io2_oeb 5.09fF
C11813 raven_soc_0|ram_wenb raven_soc_0|ram_wdata<12> 3.91fF
C11814 raven_spi_0|sdo_enb raven_soc_0|flash_io3_oeb 0.57fF
C11815 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<1> 10.18fF
C11816 LOGIC0_3V_4|Q raven_padframe_0|BBCUD4F_13|PO 0.04fF
C11817 BU_3VX2_7|A BU_3VX2_16|A 1.27fF
C11818 BU_3VX2_7|A BU_3VX2_29|A 0.01fF
C11819 LS_3VX2_7|Q LS_3VX2_6|Q 4.15fF
C11820 BU_3VX2_32|A BU_3VX2_64|A 0.52fF
C11821 BU_3VX2_6|A BU_3VX2_27|A 0.01fF
C11822 BU_3VX2_21|A raven_soc_0|flash_clk 1.72fF
C11823 raven_soc_0|gpio_pullup<1> raven_soc_0|gpio_outenb<9> 0.01fF
C11824 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<13> 4.50fF
C11825 raven_padframe_0|BBCUD4F_11|VDDR raven_padframe_0|BBCUD4F_11|VDDO 0.06fF
C11826 raven_soc_0|gpio_in<4> raven_padframe_0|BBCUD4F_4|PO 0.04fF
C11827 BU_3VX2_73|Q BU_3VX2_43|Q 0.03fF
C11828 raven_soc_0|ram_wdata<9> vdd 0.56fF
C11829 raven_soc_0|ram_wdata<1> vdd 0.38fF
C11830 BU_3VX2_54|A BU_3VX2_54|Q 0.10fF
C11831 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pullup<10> 0.01fF
C11832 BU_3VX2_9|A BU_3VX2_21|A 1.04fF
C11833 BU_3VX2_7|A BU_3VX2_37|A 1.34fF
C11834 vdd raven_padframe_0|VDDPADF_0|GNDO 0.07fF
C11835 LS_3VX2_8|Q LS_3VX2_7|Q 5.11fF
C11836 LS_3VX2_10|A LS_3VX2_9|Q 0.16fF
C11837 BU_3VX2_22|A BU_3VX2_28|A 3.65fF
C11838 raven_soc_0|gpio_out<0> raven_soc_0|gpio_pulldown<5> 0.10fF
C11839 BU_3VX2_31|A BU_3VX2_14|A 0.01fF
C11840 IN_3VX2_1|A raven_soc_0|gpio_pullup<12> 0.01fF
C11841 raven_soc_0|gpio_in<3> BU_3VX2_0|Q 0.14fF
C11842 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_outenb<7> 4.03fF
C11843 raven_soc_0|gpio_pullup<10> raven_soc_0|gpio_outenb<5> 0.47fF
C11844 raven_soc_0|gpio_pullup<9> raven_soc_0|gpio_outenb<6> 0.29fF
C11845 BU_3VX2_0|Q raven_soc_0|gpio_out<9> 0.01fF
C11846 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_out<5> 0.01fF
C11847 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_outenb<10> 3.30fF
C11848 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_out<12> 0.02fF
C11849 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<5> 0.60fF
C11850 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<6> 61.23fF
C11851 raven_soc_0|ram_wdata<6> raven_soc_0|ram_wdata<0> 4.06fF
C11852 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<15> 0.04fF
C11853 raven_soc_0|ram_rdata<8> raven_soc_0|ram_wdata<8> 0.35fF
C11854 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<8> 0.02fF
C11855 raven_soc_0|ram_rdata<5> raven_soc_0|ram_wdata<13> 0.26fF
C11856 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<6> 0.06fF
C11857 raven_soc_0|flash_io3_do raven_soc_0|flash_io2_do 322.70fF
C11858 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<1> 0.07fF
C11859 raven_soc_0|ram_rdata<9> raven_soc_0|ram_rdata<12> 14.55fF
C11860 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<14> 0.02fF
C11861 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<7> 1.80fF
C11862 raven_soc_0|ram_rdata<18> raven_soc_0|ram_wdata<14> 1.17fF
C11863 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<18> 0.27fF
C11864 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<17> 0.08fF
C11865 BU_3VX2_6|Q BU_3VX2_14|Q 4.29fF
C11866 raven_soc_0|ram_wdata<16> raven_soc_0|ram_addr<3> 0.01fF
C11867 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<4> 3.01fF
C11868 raven_soc_0|ram_wdata<10> raven_soc_0|ram_rdata<2> 0.01fF
C11869 BU_3VX2_14|Q BU_3VX2_7|Q 5.63fF
C11870 BU_3VX2_70|Q BU_3VX2_65|Q 17.02fF
C11871 LS_3VX2_23|A AMUX4_3V_3|SEL[0] 14.14fF
C11872 BU_3VX2_32|Q BU_3VX2_64|Q 3.60fF
C11873 AMUX4_3V_4|AIN2 BU_3VX2_62|Q 0.01fF
C11874 BU_3VX2_26|Q BU_3VX2_24|Q 131.85fF
C11875 vdd BU_3VX2_72|Q 2.78fF
C11876 VDD3V3 raven_padframe_0|VDDORPADF_0|GNDO 2.41fF
C11877 raven_spi_0|CSB raven_soc_0|gpio_outenb<15> 2.13fF
C11878 LOGIC0_3V_4|Q raven_soc_0|gpio_outenb<14> 10.59fF
C11879 raven_padframe_0|aregc01_3v3_0|VDDR raven_padframe_0|aregc01_3v3_0|VDDO 0.04fF
C11880 raven_padframe_0|BBCUD4F_2|GNDR raven_padframe_0|BBCUD4F_2|GNDO 0.81fF
C11881 raven_spi_0|SDO raven_soc_0|gpio_out<15> 1.97fF
C11882 AMUX4_3V_1|AIN1 LS_3VX2_17|Q 1.36fF
C11883 IN_3VX2_1|Q BU_3VX2_57|Q 0.01fF
C11884 VDD raven_padframe_0|BBCUD4F_3|GNDR 0.16fF
C11885 LS_3VX2_4|A LS_3VX2_17|A 1.18fF
C11886 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<27> 0.02fF
C11887 raven_soc_0|ram_rdata<28> raven_soc_0|ram_rdata<17> 6.22fF
C11888 LS_3VX2_19|A BU_3VX2_59|Q 12.58fF
C11889 BU_3VX2_59|Q BU_3VX2_52|Q 19.50fF
C11890 LS_3VX2_12|A VDD3V3 0.51fF
C11891 BU_3VX2_35|A raven_soc_0|ext_clk 0.17fF
C11892 LS_3VX2_14|A LS_3VX2_27|A 11.66fF
C11893 BU_3VX2_65|A BU_3VX2_66|Q 0.03fF
C11894 BU_3VX2_69|A BU_3VX2_67|Q 0.03fF
C11895 BU_3VX2_0|Q raven_soc_0|ram_rdata<21> 0.02fF
C11896 BU_3VX2_26|A raven_soc_0|flash_io0_di 0.01fF
C11897 BU_3VX2_31|A apllc03_1v8_0|B_CP 5.26fF
C11898 BU_3VX2_63|Q raven_soc_0|gpio_in<8> 0.01fF
C11899 raven_soc_0|gpio_pulldown<1> BU_3VX2_29|Q 0.01fF
C11900 raven_soc_0|gpio_pulldown<15> raven_soc_0|ext_clk 0.01fF
C11901 IN_3VX2_1|A BU_3VX2_53|Q 0.01fF
C11902 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_in<13> 10.13fF
C11903 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_in<9> 0.01fF
C11904 raven_soc_0|gpio_in<2> BU_3VX2_72|Q 0.13fF
C11905 BU_3VX2_27|A BU_3VX2_25|Q 0.03fF
C11906 BU_3VX2_7|A LS_3VX2_3|Q 0.98fF
C11907 BU_3VX2_32|A BU_3VX2_66|A 0.54fF
C11908 raven_padframe_0|FILLER20F_0|VDDR raven_padframe_0|FILLER20F_0|VDDO 0.06fF
C11909 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_pulldown<12> 0.01fF
C11910 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_outenb<0> 29.63fF
C11911 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<4> 0.01fF
C11912 BU_3VX2_11|A raven_soc_0|flash_io0_di 0.01fF
C11913 raven_soc_0|gpio_in<3> raven_soc_0|flash_io3_di 0.28fF
C11914 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pulldown<7> 13.18fF
C11915 BU_3VX2_63|Q raven_soc_0|gpio_pullup<13> 0.09fF
C11916 adc_low BU_3VX2_59|Q 0.05fF
C11917 raven_padframe_0|FILLER20F_5|VDDR raven_padframe_0|FILLER20F_5|VDDO 0.06fF
C11918 raven_soc_0|gpio_in<6> raven_soc_0|irq_pin 0.01fF
C11919 BU_3VX2_73|Q BU_3VX2_50|Q 12.80fF
C11920 raven_padframe_0|BT4FC_0|VDDR raven_padframe_0|BT4FC_0|VDD3 0.71fF
C11921 BU_3VX2_3|A BU_3VX2_19|A 0.01fF
C11922 BU_3VX2_19|A BU_3VX2_15|A 4.98fF
C11923 BU_3VX2_21|A BU_3VX2_28|A 3.04fF
C11924 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pulldown<13> 0.01fF
C11925 BU_3VX2_38|A raven_soc_0|flash_csb 0.01fF
C11926 LS_3VX2_4|Q LS_3VX2_24|Q 0.01fF
C11927 raven_soc_0|ram_addr<5> raven_soc_0|ram_addr<9> 10.94fF
C11928 raven_soc_0|ram_addr<6> raven_soc_0|ram_addr<8> 30.74fF
C11929 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<15> 0.11fF
C11930 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<13> 0.40fF
C11931 raven_soc_0|ram_wdata<19> raven_soc_0|ram_wdata<29> 7.95fF
C11932 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<13> 4.56fF
C11933 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<0> 0.10fF
C11934 raven_soc_0|ram_addr<9> raven_soc_0|ram_wdata<19> 0.01fF
C11935 raven_soc_0|ram_rdata<29> raven_soc_0|ram_wdata<31> 0.01fF
C11936 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<16> 0.01fF
C11937 raven_soc_0|ram_addr<7> raven_soc_0|ram_wdata<25> 0.01fF
C11938 raven_soc_0|ram_addr<5> raven_soc_0|ram_wdata<29> 0.01fF
C11939 raven_soc_0|ram_addr<6> raven_soc_0|ram_wdata<22> 0.01fF
C11940 BU_3VX2_56|Q LS_3VX2_27|A 0.74fF
C11941 raven_soc_0|gpio_in<15> apllc03_1v8_0|CLK 0.02fF
C11942 AMUX4_3V_1|SEL[0] vdd 3.59fF
C11943 BU_3VX2_50|A BU_3VX2_44|A 0.41fF
C11944 BU_3VX2_51|A LS_3VX2_20|Q 0.13fF
C11945 raven_soc_0|gpio_in<10> BU_3VX2_23|Q 0.01fF
C11946 raven_soc_0|gpio_out<15> BU_3VX2_26|Q 0.01fF
C11947 raven_padframe_0|VDDPADF_1|GNDR raven_padframe_0|VDDPADF_1|VDDO 0.09fF
C11948 BU_3VX2_22|A BU_3VX2_14|A 2.08fF
C11949 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_pullup<1> 13.31fF
C11950 raven_padframe_0|aregc01_3v3_1|m4_92500_28769# raven_padframe_0|aregc01_3v3_1|m4_92500_22024# 0.03fF
C11951 BU_3VX2_63|Q raven_soc_0|gpio_out<5> 0.01fF
C11952 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_outenb<10> 0.01fF
C11953 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<14> 0.67fF
C11954 LS_3VX2_10|A BU_3VX2_73|Q 7.89fF
C11955 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<10> 3.68fF
C11956 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<5> 27.56fF
C11957 BU_3VX2_0|Q raven_soc_0|ext_clk 27.49fF
C11958 raven_soc_0|gpio_pulldown<10> raven_soc_0|gpio_in<9> 9.91fF
C11959 raven_soc_0|gpio_pulldown<9> VDD3V3 0.07fF
C11960 BU_3VX2_71|Q vdd 1.03fF
C11961 raven_soc_0|gpio_outenb<13> BU_3VX2_24|Q 0.01fF
C11962 raven_soc_0|gpio_pullup<14> BU_3VX2_28|Q 0.01fF
C11963 BU_3VX2_36|Q vdd 1.28fF
C11964 BU_3VX2_37|Q BU_3VX2_27|Q 0.02fF
C11965 BU_3VX2_11|Q BU_3VX2_24|Q 2.81fF
C11966 BU_3VX2_8|A raven_soc_0|flash_io2_do 0.01fF
C11967 BU_3VX2_7|A raven_soc_0|flash_io1_oeb 0.01fF
C11968 IN_3VX2_1|Q LS_3VX2_16|A 0.01fF
C11969 LS_3VX2_2|Q vdd 0.12fF
C11970 raven_padframe_0|VDDPADF_1|VDDR raven_padframe_0|VDDPADF_1|GNDO 0.13fF
C11971 BU_3VX2_17|A BU_3VX2_15|Q 0.03fF
C11972 BU_3VX2_18|A raven_soc_0|flash_io3_oeb 0.01fF
C11973 BU_3VX2_31|A raven_soc_0|flash_io1_do 5.98fF
C11974 raven_soc_0|gpio_pulldown<0> raven_soc_0|ext_clk 0.01fF
C11975 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pulldown<3> 2.68fF
C11976 raven_soc_0|gpio_in<3> raven_soc_0|irq_pin 0.01fF
C11977 LS_3VX2_3|A raven_soc_0|gpio_out<8> 0.86fF
C11978 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_pullup<14> 10.16fF
C11979 BU_3VX2_0|Q raven_soc_0|ram_rdata<17> 0.02fF
C11980 raven_soc_0|ram_rdata<20> raven_soc_0|ram_rdata<23> 29.86fF
C11981 raven_soc_0|ram_rdata<0> raven_soc_0|ram_rdata<19> 0.79fF
C11982 BU_3VX2_48|A BU_3VX2_45|A 0.92fF
C11983 BU_3VX2_59|Q BU_3VX2_58|Q 237.81fF
C11984 BU_3VX2_48|A BU_3VX2_47|Q 0.15fF
C11985 raven_padframe_0|APR00DF_6|VDDO raven_padframe_0|APR00DF_6|GNDO 2.28fF
C11986 LS_3VX2_6|Q LS_3VX2_4|Q 0.96fF
C11987 BU_3VX2_23|A raven_soc_0|flash_io0_do 0.01fF
C11988 BU_3VX2_40|A BU_3VX2_71|Q 0.03fF
C11989 raven_soc_0|gpio_out<0> BU_3VX2_29|Q 0.01fF
C11990 raven_padframe_0|ICFC_1|VDDR raven_padframe_0|ICFC_1|GNDO 0.13fF
C11991 raven_soc_0|gpio_in<2> BU_3VX2_71|Q 0.14fF
C11992 BU_3VX2_13|A BU_3VX2_11|Q 0.03fF
C11993 raven_soc_0|gpio_out<2> raven_soc_0|gpio_pullup<13> 0.08fF
C11994 BU_3VX2_33|A BU_3VX2_32|Q 0.16fF
C11995 raven_soc_0|gpio_in<0> BU_3VX2_23|Q 0.01fF
C11996 LOGIC0_3V_4|Q raven_padframe_0|ICF_0|PO 0.04fF
C11997 AMUX2_3V_0|SEL BU_3VX2_52|Q 0.01fF
C11998 raven_soc_0|gpio_out<12> BU_3VX2_29|Q 0.01fF
C11999 raven_soc_0|flash_csb BU_3VX2_23|Q 0.01fF
C12000 raven_soc_0|gpio_out<13> apllc03_1v8_0|CLK 0.01fF
C12001 BU_3VX2_54|A BU_3VX2_56|Q 0.04fF
C12002 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<4> 0.01fF
C12003 LS_3VX2_8|Q LS_3VX2_4|Q 0.45fF
C12004 VDD raven_soc_0|gpio_pullup<15> 0.27fF
C12005 BU_3VX2_5|A BU_3VX2_26|A 0.01fF
C12006 LS_3VX2_5|Q LS_3VX2_6|A 0.16fF
C12007 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<0> 0.01fF
C12008 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<14> 0.01fF
C12009 IN_3VX2_1|A raven_soc_0|gpio_outenb<0> 0.01fF
C12010 raven_soc_0|gpio_outenb<1> raven_soc_0|gpio_pulldown<11> 0.01fF
C12011 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_outenb<14> 45.99fF
C12012 raven_soc_0|gpio_pullup<8> raven_soc_0|gpio_pullup<9> 15.90fF
C12013 raven_soc_0|gpio_pullup<3> raven_soc_0|gpio_pullup<12> 0.01fF
C12014 raven_soc_0|gpio_pullup<4> raven_soc_0|gpio_pullup<11> 0.18fF
C12015 raven_soc_0|gpio_pullup<7> raven_soc_0|gpio_pullup<10> 1.27fF
C12016 LS_3VX2_3|A raven_soc_0|gpio_out<6> 0.01fF
C12017 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_outenb<6> 0.01fF
C12018 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_outenb<12> 0.02fF
C12019 BU_3VX2_0|Q raven_soc_0|gpio_outenb<10> 0.01fF
C12020 raven_soc_0|ram_wdata<4> raven_soc_0|ram_wdata<6> 21.22fF
C12021 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<31> 0.02fF
C12022 raven_soc_0|ram_wdata<9> raven_soc_0|ram_rdata<24> 2.01fF
C12023 raven_soc_0|ram_wdata<5> raven_soc_0|ram_wdata<23> 0.01fF
C12024 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<10> 8.75fF
C12025 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<5> 0.01fF
C12026 raven_soc_0|ram_rdata<24> raven_soc_0|ram_wdata<1> 2.07fF
C12027 raven_soc_0|ram_wdata<10> raven_soc_0|ram_wdata<2> 4.53fF
C12028 raven_soc_0|ram_rdata<14> raven_soc_0|ram_rdata<12> 28.01fF
C12029 AMUX4_3V_3|SEL[1] BU_3VX2_22|Q 0.45fF
C12030 raven_soc_0|ram_rdata<22> raven_soc_0|ram_wdata<8> 0.28fF
C12031 raven_soc_0|ram_wdata<23> raven_soc_0|ram_wdata<0> 0.01fF
C12032 raven_soc_0|ext_clk raven_soc_0|flash_io3_di 42.37fF
C12033 raven_soc_0|flash_io0_di VDD3V3 9.23fF
C12034 LS_3VX2_17|A vdd 1.09fF
C12035 VDD3V3 BU_3VX2_46|Q 0.24fF
C12036 vdd apllc03_1v8_0|VCO_IN 0.04fF
C12037 BU_3VX2_21|A BU_3VX2_14|A 2.43fF
C12038 BU_3VX2_5|A BU_3VX2_11|A 1.82fF
C12039 LOGIC0_3V_4|Q raven_soc_0|gpio_pullup<15> 107.05fF
C12040 raven_padframe_0|aregc01_3v3_0|m4_92500_30133# raven_padframe_0|aregc01_3v3_0|GNDR 0.07fF
C12041 adc_low AMUX2_3V_0|SEL 0.05fF
C12042 raven_soc_0|gpio_out<2> raven_soc_0|gpio_out<5> 0.46fF
C12043 AMUX4_3V_1|AIN1 BU_3VX2_54|A 0.02fF
C12044 BU_3VX2_12|A BU_3VX2_9|Q 0.02fF
C12045 raven_soc_0|ram_addr<1> raven_soc_0|ram_rdata<19> 0.32fF
C12046 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<21> 0.03fF
C12047 BU_3VX2_71|Q raven_soc_0|gpio_in<11> 0.41fF
C12048 raven_soc_0|ram_rdata<19> raven_soc_0|ram_wdata<26> 0.01fF
C12049 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<15> 0.02fF
C12050 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_out<15> 12.45fF
C12051 raven_soc_0|ram_addr<8> raven_soc_0|ram_rdata<28> 4.06fF
C12052 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<25> 0.01fF
C12053 LS_3VX2_22|A BU_3VX2_59|Q 0.03fF
C12054 raven_soc_0|ram_wdata<6> vdd 0.55fF
C12055 LS_3VX2_19|A BU_3VX2_61|Q 19.26fF
C12056 BU_3VX2_61|Q BU_3VX2_52|Q 13.95fF
C12057 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pulldown<1> 24.77fF
C12058 BU_3VX2_24|A BU_3VX2_22|Q 0.03fF
C12059 LS_3VX2_8|A BU_3VX2_42|Q 6.21fF
C12060 raven_soc_0|gpio_outenb<3> vdd 0.37fF
C12061 raven_soc_0|gpio_outenb<9> BU_3VX2_71|Q 0.49fF
C12062 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<5> 0.01fF
C12063 raven_soc_0|ram_rdata<6> raven_soc_0|ram_wdata<6> 0.44fF
C12064 raven_soc_0|ram_addr<2> raven_soc_0|ram_rdata<31> 21.32fF
C12065 raven_soc_0|ram_rdata<9> raven_soc_0|ram_wdata<24> 0.02fF
C12066 raven_soc_0|ram_wdata<20> raven_soc_0|ram_rdata<10> 0.33fF
C12067 BU_3VX2_70|Q BU_3VX2_36|Q 1.32fF
C12068 raven_padframe_0|BBC4F_2|VDDO raven_padframe_0|BBC4F_2|GNDO 2.28fF
C12069 raven_padframe_0|BBCUD4F_14|VDDO raven_padframe_0|BBCUD4F_14|GNDO 2.28fF
C12070 raven_padframe_0|BBCUD4F_8|VDDO raven_padframe_0|BBCUD4F_8|GNDO 2.28fF
C12071 markings_0|manufacturer_0|_alphabet_B_0|m2_0_0# markings_0|product_name_0|_alphabet_E_0|m2_0_0# 0.35fF
C12072 raven_soc_0|gpio_in<1> raven_soc_0|flash_io2_di 0.26fF
C12073 BU_3VX2_22|A raven_soc_0|flash_io1_do 0.01fF
C12074 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<10> 0.01fF
C12075 raven_soc_0|gpio_pulldown<2> LS_3VX2_3|A 0.01fF
C12076 LS_3VX2_23|Q vdd 1.66fF
C12077 BU_3VX2_71|A raven_soc_0|flash_io3_oeb 0.01fF
C12078 IN_3VX2_1|A raven_soc_0|flash_io0_do 5.93fF
C12079 raven_soc_0|gpio_outenb<4> raven_soc_0|gpio_pullup<6> 0.23fF
C12080 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pulldown<3> 0.46fF
C12081 VDD raven_padframe_0|BBCUD4F_11|GNDO 0.07fF
C12082 adc_low BU_3VX2_61|Q 0.05fF
C12083 raven_soc_0|ext_clk raven_soc_0|irq_pin 0.07fF
C12084 BU_3VX2_73|Q BU_3VX2_48|Q 9.67fF
C12085 BU_3VX2_2|A BU_3VX2_71|A 0.01fF
C12086 LS_3VX2_7|Q LS_3VX2_14|Q 0.40fF
C12087 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_in<2> 6.47fF
C12088 raven_soc_0|gpio_out<11> raven_soc_0|gpio_out<14> 1.30fF
C12089 raven_soc_0|gpio_out<13> raven_soc_0|gpio_outenb<8> 1.90fF
C12090 AMUX2_3V_0|SEL BU_3VX2_58|Q 0.01fF
C12091 raven_soc_0|ram_rdata<26> raven_soc_0|ram_addr<7> 3.86fF
C12092 raven_soc_0|ram_rdata<27> raven_soc_0|ram_addr<6> 4.37fF
C12093 raven_soc_0|ram_wdata<30> raven_soc_0|ram_addr<9> 0.01fF
C12094 raven_soc_0|ram_rdata<29> raven_soc_0|ram_addr<5> 6.25fF
C12095 raven_soc_0|ram_wdata<12> raven_soc_0|ram_rdata<13> 0.05fF
C12096 BU_3VX2_21|Q BU_3VX2_17|Q 8.99fF
C12097 raven_soc_0|ram_wdata<30> raven_soc_0|ram_wdata<29> 188.12fF
C12098 raven_soc_0|ram_wdata<17> raven_soc_0|ram_wdata<21> 21.99fF
C12099 raven_soc_0|ram_rdata<2> raven_soc_0|ram_wdata<25> 2.10fF
C12100 raven_soc_0|ram_rdata<25> raven_soc_0|ram_wdata<31> 0.10fF
C12101 BU_3VX2_73|Q raven_soc_0|ser_tx 0.01fF
C12102 BU_3VX2_1|Q BU_3VX2_69|Q 0.54fF
C12103 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<27> 4.55fF
C12104 raven_soc_0|gpio_in<13> BU_3VX2_23|Q 0.01fF
C12105 BU_3VX2_8|Q BU_3VX2_17|Q 7.39fF
C12106 AMUX4_3V_4|AIN3 AMUX4_3V_4|AIN2 55.98fF
C12107 raven_soc_0|gpio_in<14> apllc03_1v8_0|CLK 0.13fF
C12108 BU_3VX2_33|Q BU_3VX2_52|Q 0.39fF
C12109 raven_soc_0|gpio_in<9> BU_3VX2_28|Q 0.01fF
C12110 BU_3VX2_40|Q BU_3VX2_27|Q 2.00fF
C12111 BU_3VX2_54|Q BU_3VX2_53|Q 231.64fF
C12112 raven_soc_0|gpio_in<1> raven_soc_0|gpio_pulldown<11> 0.01fF
C12113 LS_3VX2_9|A LS_3VX2_13|A 10.39fF
C12114 raven_padframe_0|aregc01_3v3_1|m4_92500_30653# raven_padframe_0|aregc01_3v3_1|m4_92500_30133# 0.09fF
C12115 raven_padframe_0|aregc01_3v3_1|m4_92500_31172# raven_padframe_0|aregc01_3v3_1|m4_92500_29333# 0.01fF
C12116 IN_3VX2_1|A raven_soc_0|gpio_pulldown<14> 0.01fF
C12117 raven_soc_0|gpio_pulldown<8> raven_soc_0|gpio_pullup<4> 0.12fF
C12118 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pullup<10> 0.01fF
C12119 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_outenb<5> 0.01fF
C12120 BU_3VX2_63|Q raven_soc_0|gpio_outenb<6> 0.01fF
C12121 BU_3VX2_63|A raven_soc_0|ext_clk 0.01fF
C12122 LS_3VX2_24|A BU_3VX2_73|Q 164.77fF
C12123 raven_soc_0|gpio_out<4> raven_soc_0|gpio_in<13> 0.02fF
C12124 raven_soc_0|gpio_pulldown<12> raven_soc_0|gpio_in<9> 0.01fF
C12125 BU_3VX2_1|Q raven_soc_0|flash_io0_oeb 0.66fF
C12126 raven_soc_0|gpio_pullup<14> vdd 0.37fF
C12127 raven_soc_0|gpio_out<10> BU_3VX2_26|Q 0.01fF
C12128 raven_soc_0|gpio_pullup<13> BU_3VX2_24|Q 0.01fF
C12129 raven_soc_0|gpio_pullup<6> apllc03_1v8_0|CLK 0.01fF
C12130 BU_3VX2_37|Q BU_3VX2_25|Q 0.53fF
C12131 BU_3VX2_14|Q BU_3VX2_23|Q 10.15fF
C12132 LOGIC0_3V_4|Q raven_soc_0|gpio_out<3> 0.01fF
C12133 BU_3VX2_5|A VDD3V3 0.24fF
C12134 BU_3VX2_19|A BU_3VX2_17|Q 0.03fF
C12135 BU_3VX2_31|A raven_soc_0|gpio_in<10> 0.01fF
C12136 VDD raven_padframe_0|GNDORPADF_2|VDDR 0.71fF
C12137 raven_spi_0|sdo_enb raven_soc_0|gpio_in<15> 1.32fF
C12138 LS_3VX2_3|A raven_soc_0|gpio_pulldown<6> 0.14fF
C12139 raven_soc_0|gpio_out<2> VDD3V3 2.25fF
C12140 BU_3VX2_0|Q raven_soc_0|ram_wdata<22> 0.02fF
C12141 BU_3VX2_26|A BU_3VX2_24|Q 0.03fF
C12142 raven_soc_0|ser_rx raven_padframe_0|ICF_0|PO 0.04fF
C12143 BU_3VX2_51|A BU_3VX2_47|A 1.39fF
C12144 BU_3VX2_50|A BU_3VX2_48|A 4.05fF
C12145 BU_3VX2_61|Q BU_3VX2_58|Q 49.13fF
C12146 BU_3VX2_60|Q BU_3VX2_59|Q 232.36fF
C12147 BU_3VX2_49|A adc0_data<5> 0.02fF
C12148 raven_padframe_0|VDDORPADF_0|GNDR raven_padframe_0|VDDORPADF_0|GNDO 0.81fF
C12149 raven_padframe_0|APR00DF_6|VDDR raven_padframe_0|APR00DF_6|VDDO 0.06fF
C12150 raven_soc_0|gpio_out<1> raven_soc_0|gpio_out<0> 18.03fF
C12151 raven_padframe_0|APR00DF_4|VDDR raven_padframe_0|APR00DF_4|VDDO 0.06fF
C12152 BU_3VX2_73|A adc_high 0.09fF
C12153 BU_3VX2_23|A raven_soc_0|flash_io1_di 0.01fF
C12154 BU_3VX2_21|A raven_soc_0|flash_io1_do 0.01fF
C12155 raven_soc_0|gpio_outenb<3> raven_soc_0|gpio_outenb<9> 0.77fF
C12156 VDD raven_padframe_0|APR00DF_6|GNDR 0.16fF
C12157 raven_soc_0|gpio_in<2> raven_soc_0|gpio_pullup<14> 0.01fF
C12158 raven_soc_0|gpio_outenb<2> raven_soc_0|gpio_pulldown<7> 0.01fF
C12159 AMUX2_3V_0|SEL LS_3VX2_22|A 170.86fF
C12160 raven_padframe_0|BBCUD4F_8|VDDR raven_padframe_0|BBCUD4F_8|GNDO 0.13fF
C12161 raven_soc_0|gpio_outenb<12> BU_3VX2_29|Q 0.01fF
C12162 raven_soc_0|gpio_outenb<15> apllc03_1v8_0|CLK 0.01fF
C12163 raven_padframe_0|BBCUD4F_4|VDDR raven_padframe_0|BBCUD4F_4|GNDO 0.13fF
C12164 BU_3VX2_33|A raven_padframe_0|ICFC_2|PO 0.04fF
C12165 raven_soc_0|gpio_out<9> BU_3VX2_26|Q 0.01fF
C12166 LS_3VX2_9|A raven_soc_0|ser_rx 0.01fF
C12167 BU_3VX2_66|A BU_3VX2_64|A 8.38fF
C12168 BU_3VX2_13|A BU_3VX2_26|A 1.61fF
C12169 raven_soc_0|gpio_pullup<2> BU_3VX2_71|Q 0.01fF
C12170 IN_3VX2_1|A raven_soc_0|gpio_pulldown<10> 0.01fF
C12171 raven_soc_0|gpio_pulldown<4> raven_soc_0|gpio_pullup<7> 0.03fF
C12172 LS_3VX2_3|A raven_soc_0|gpio_outenb<11> 0.01fF
C12173 BU_3VX2_0|Q raven_soc_0|gpio_pullup<10> 0.01fF
C12174 raven_soc_0|gpio_pulldown<13> raven_soc_0|gpio_pullup<15> 11.41fF
C12175 raven_soc_0|gpio_pulldown<5> raven_soc_0|gpio_pullup<12> 0.02fF
C12176 BU_3VX2_25|A raven_soc_0|flash_io0_do 2.50fF
C12177 raven_soc_0|gpio_outenb<0> raven_soc_0|gpio_pullup<3> 0.01fF
C12178 raven_soc_0|gpio_pulldown<9> raven_soc_0|gpio_pullup<8> 15.44fF
C12179 raven_soc_0|ram_wdata<3> raven_soc_0|ram_rdata<30> 0.11fF
C12180 raven_soc_0|ram_wenb raven_soc_0|ram_addr<4> 0.01fF
C12181 AMUX4_3V_3|SEL[1] BU_3VX2_31|Q 1.64fF
C12182 BU_3VX2_40|Q raven_soc_0|flash_io2_oeb 0.02fF
C12183 raven_soc_0|gpio_in<8> raven_soc_0|gpio_out<15> 0.01fF
C12184 BU_3VX2_42|Q BU_3VX2_44|Q 28.86fF
C12185 AMUX4_3V_0|SEL[1] BU_3VX2_51|Q 9.12fF
C12186 BU_3VX2_13|A BU_3VX2_11|A 13.03fF
C12187 BU_3VX2_31|A raven_soc_0|gpio_in<0> 0.01fF
C12188 raven_padframe_0|aregc01_3v3_0|m4_92500_30653# raven_padframe_0|aregc01_3v3_0|m4_92500_29333# 0.02fF
C12189 raven_padframe_0|aregc01_3v3_0|m4_0_29057# raven_padframe_0|aregc01_3v3_0|m4_0_22024# 0.02fF
C12190 BU_3VX2_31|A raven_soc_0|flash_csb 165.43fF
C12191 raven_soc_0|gpio_out<2> raven_soc_0|gpio_outenb<6> 0.01fF
C12192 raven_soc_0|gpio_outenb<8> raven_soc_0|gpio_in<14> 0.02fF
C12193 raven_soc_0|ram_rdata<27> raven_soc_0|ram_rdata<28> 168.95fF
C12194 raven_soc_0|gpio_out<14> raven_soc_0|gpio_in<12> 14.39fF
C12195 raven_soc_0|ram_rdata<3> raven_soc_0|ram_rdata<20> 2.48fF
C12196 raven_soc_0|gpio_in<5> raven_soc_0|gpio_in<8> 1.14fF
C12197 raven_soc_0|ram_wdata<18> raven_soc_0|ram_rdata<23> 0.25fF
C12198 raven_soc_0|gpio_out<8> raven_soc_0|gpio_in<10> 3.40fF
C12199 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<11> 0.01fF
C12200 raven_soc_0|gpio_outenb<13> raven_soc_0|gpio_in<6> 0.01fF
C12201 raven_soc_0|gpio_pullup<14> raven_soc_0|gpio_in<11> 0.01fF
C12202 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_out<15> 20.64fF
C12203 raven_soc_0|ram_wdata<28> raven_soc_0|ram_rdata<19> 0.01fF
C12204 raven_soc_0|ram_rdata<0> raven_soc_0|ram_wdata<15> 0.17fF
C12205 raven_soc_0|ram_rdata<11> raven_soc_0|ram_wdata<13> 0.02fF
C12206 raven_soc_0|ram_rdata<20> raven_soc_0|ram_wdata<14> 0.01fF
C12207 LS_3VX2_22|A BU_3VX2_61|Q 0.12fF
C12208 raven_soc_0|ram_wdata<23> vdd 0.66fF
C12209 LS_3VX2_19|A LS_3VX2_15|A 23.34fF
C12210 LS_3VX2_15|A BU_3VX2_52|Q 9.50fF
C12211 raven_spi_0|CSB LOGIC0_3V_4|Q 0.94fF
C12212 raven_soc_0|gpio_in<5> raven_padframe_0|BBCUD4F_5|PO 0.04fF
C12213 VDD raven_padframe_0|BBC4F_1|GNDR 0.16fF
C12214 LS_3VX2_14|A BU_3VX2_53|Q 0.02fF
C12215 raven_soc_0|gpio_pullup<0> BU_3VX2_28|Q 0.01fF
C12216 raven_soc_0|gpio_outenb<1> BU_3VX2_23|Q 0.01fF
C12217 raven_soc_0|gpio_pullup<6> raven_soc_0|gpio_outenb<8> 6.73fF
C12218 raven_soc_0|gpio_outenb<9> raven_soc_0|gpio_pullup<14> 1.14fF
C12219 raven_soc_0|gpio_out<10> raven_soc_0|gpio_outenb<13> 0.26fF
C12220 raven_soc_0|gpio_pullup<13> raven_soc_0|gpio_in<5> 0.01fF
C12221 raven_soc_0|ram_rdata<18> raven_soc_0|ram_rdata<31> 6.13fF
C12222 raven_soc_0|ram_rdata<21> raven_soc_0|ram_rdata<10> 3.47fF
C12223 raven_soc_0|ram_rdata<30> raven_soc_0|ram_addr<2> 15.48fF
C12224 raven_soc_0|ram_rdata<8> raven_soc_0|ram_rdata<9> 64.58fF
C12225 raven_soc_0|ram_wdata<23> raven_soc_0|ram_rdata<6> 0.67fF
C12226 BU_3VX2_14|Q BU_3VX2_4|Q 5.95fF
C12227 raven_soc_0|ram_rdata<14> raven_soc_0|ram_wdata<24> 0.02fF
C12228 raven_soc_0|ram_addr<3> raven_soc_0|ram_wdata<20> 0.01fF
C12229 raven_soc_0|ram_rdata<4> raven_soc_0|ram_wdata<7> 0.01fF
C12230 BU_3VX2_24|A raven_soc_0|flash_io3_oeb 2.75fF
C12231 BU_3VX2_3|A raven_soc_0|flash_io2_oeb 0.01fF
C12232 raven_soc_0|gpio_pullup<0> raven_soc_0|gpio_pulldown<12> 0.01fF
C12233 AMUX4_3V_3|AOUT AMUX4_3V_4|AIN3 23.67fF
C12234 BU_3VX2_15|A raven_soc_0|flash_io2_oeb 0.01fF
C12235 raven_padframe_0|BBC4F_0|VDDR raven_padframe_0|BBC4F_0|GNDR 0.68fF
C12236 IN_3VX2_1|A raven_soc_0|flash_io1_di 0.01fF
C12237 adc_low LS_3VX2_15|A 0.05fF
C12238 raven_soc_0|gpio_out<13> raven_soc_0|gpio_in<15> 12.65fF
C12239 raven_soc_0|gpio_out<6> raven_soc_0|gpio_in<10> 0.49fF
C12240 VDD raven_padframe_0|BBCUD4F_4|GNDR 0.16fF
C12241 BU_3VX2_24|A BU_3VX2_2|A 0.01fF
C12242 BU_3VX2_23|A BU_3VX2_10|A 0.96fF
C12243 BU_3VX2_3|A BU_3VX2_6|A 4.36fF
C12244 BU_3VX2_6|A BU_3VX2_15|A 1.23fF
C12245 BU_3VX2_20|A BU_3VX2_31|A 1.91fF
C12246 LS_3VX2_4|Q LS_3VX2_14|Q 5.27fF
C12247 AMUX4_3V_0|AIN1 BU_3VX2_49|A 0.02fF
C12248 raven_soc_0|gpio_in<0> raven_soc_0|gpio_out<8> 0.05fF
C12249 raven_soc_0|gpio_out<1> raven_soc_0|gpio_pullup<5> 0.01fF
C12250 raven_soc_0|gpio_in<3> raven_soc_0|gpio_outenb<13> 0.01fF
C12251 raven_soc_0|gpio_out<9> raven_soc_0|gpio_outenb<13> 0.04fF
C12252 raven_soc_0|gpio_outenb<15> raven_soc_0|gpio_outenb<8> 0.03fF
C12253 raven_soc_0|gpio_outenb<14> BU_3VX2_71|Q 0.01fF
C12254 AMUX2_3V_0|SEL BU_3VX2_60|Q 0.01fF
C12255 raven_soc_0|ram_wdata<30> raven_soc_0|ram_rdata<29> 0.13fF
C12256 BU_3VX2_15|Q BU_3VX2_2|Q 2.52fF
C12257 raven_soc_0|ram_rdata<26> raven_soc_0|ram_rdata<2> 2.75fF
C12258 BU_3VX2_12|Q BU_3VX2_13|Q 68.58fF
C12259 raven_soc_0|ram_wdata<18> raven_soc_0|ram_wdata<21> 30.94fF
C12260 raven_soc_0|ram_rdata<3> raven_soc_0|ram_wdata<17> 0.01fF
C12261 raven_soc_0|ram_addr<5> raven_soc_0|ram_rdata<25> 4.09fF
C12262 raven_soc_0|ram_wdata<16> raven_soc_0|ram_wdata<25> 8.20fF
C12263 raven_soc_0|ram_rdata<12> raven_soc_0|ram_wdata<29> 0.12fF
C12264 raven_soc_0|ram_wdata<13> raven_soc_0|ram_rdata<2> 3.01fF
C12265 BU_3VX2_18|Q BU_3VX2_17|Q 64.39fF
C12266 raven_soc_0|ram_wdata<14> raven_soc_0|ram_wdata<17> 23.13fF
C12267 BU_3VX2_2|Q BU_3VX2_9|Q 5.56fF
C12268 BU_3VX2_22|Q BU_3VX2_67|Q 20.54fF
C12269 BU_3VX2_38|Q BU_3VX2_22|Q 0.02fF
C12270 BU_3VX2_7|Q BU_3VX2_20|Q 3.30fF
C12271 BU_3VX2_19|Q BU_3VX2_17|Q 21.86fF
C12272 BU_3VX2_66|Q BU_3VX2_7|Q 0.27fF
C12273 BU_3VX2_15|Q BU_3VX2_10|Q 7.42fF
C12274 BU_3VX2_9|Q BU_3VX2_10|Q 68.48fF
C12275 raven_soc_0|ram_wdata<15> raven_soc_0|ram_wdata<26> 5.01fF
C12276 raven_soc_0|ram_wdata<8> raven_soc_0|ram_wdata<21> 2.93fF
C12277 raven_soc_0|ext_clk BU_3VX2_26|Q 0.01fF
C12278 raven_soc_0|gpio_in<9> vdd 4.45fF
C12279 BU_3VX2_40|Q BU_3VX2_25|Q 0.01fF
C12280 BU_3VX2_42|Q vdd 3.19fF
C12281 BU_3VX2_56|Q BU_3VX2_53|Q 72.39fF
C12282 BU_3VX2_57|A vdd 1.25fF
C12283 BU_3VX2_43|Q BU_3VX2_50|Q 14.57fF
C12284 VDD3V3 BU_3VX2_24|Q 0.79fF
C12285 raven_padframe_0|BBC4F_1|GNDR raven_padframe_0|BBC4F_1|VDDO 0.09fF
C12286 raven_padframe_0|FILLER50F_2|GNDR raven_padframe_0|FILLER50F_2|VDDO 0.09fF
C12287 BU_3VX2_23|A BU_3VX2_0|A 0.01fF
C12288 raven_padframe_0|FILLER20F_7|GNDR raven_padframe_0|FILLER20F_7|VDDO 0.09fF
C12289 raven_soc_0|gpio_pullup<2> raven_soc_0|gpio_outenb<3> 13.09fF
C12290 raven_padframe_0|aregc01_3v3_1|m4_0_30133# raven_padframe_0|aregc01_3v3_1|m4_0_29333# 0.09fF
C12291 raven_padframe_0|aregc01_3v3_1|m4_0_30653# raven_padframe_0|aregc01_3v3_1|m4_0_29057# 0.01fF
C12292 raven_soc_0|gpio_out<3> raven_soc_0|gpio_pulldown<13> 0.01fF
C12293 raven_padframe_0|axtoc02_3v3_0|m4_0_30653# raven_padframe_0|axtoc02_3v3_0|m4_0_30133# 0.17fF
C12294 raven_padframe_0|axtoc02_3v3_0|m4_0_31172# raven_padframe_0|axtoc02_3v3_0|m4_0_29333# 0.02fF
C12295 raven_soc_0|gpio_pulldown<14> raven_soc_0|gpio_pullup<3> 0.01fF
C12296 BU_3VX2_63|Q raven_soc_0|gpio_pullup<8> 0.01fF
C12297 raven_soc_0|gpio_pulldown<11> raven_soc_0|gpio_pullup<7> 0.01fF
C12298 raven_soc_0|gpio_pulldown<15> raven_soc_0|gpio_pulldown<4> 0.01fF
C12299 raven_padframe_0|GNDORPADF_7|VDDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12300 raven_padframe_0|GNDORPADF_1|VDDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12301 raven_padframe_0|GNDORPADF_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.81fF
C12302 raven_padframe_0|GNDORPADF_6|VDDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12303 raven_padframe_0|GNDORPADF_6|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.81fF
C12304 raven_padframe_0|GNDORPADF_2|VDDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12305 raven_padframe_0|GNDORPADF_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.81fF
C12306 raven_padframe_0|GNDORPADF_3|VDDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12307 BU_3VX2_27|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.76fF
C12308 apllc03_1v8_0|B_CP raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.91fF
C12309 BU_3VX2_29|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -19.61fF
C12310 BU_3VX2_72|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.99fF
C12311 apllc03_1v8_0|CLK raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.13fF
C12312 BU_3VX2_28|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -18.06fF
C12313 apllc03_1v8_0|B_VCO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.13fF
C12314 BU_3VX2_23|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.54fF
C12315 BU_3VX2_24|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.37fF
C12316 BU_3VX2_25|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.22fF
C12317 BU_3VX2_26|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.98fF
C12318 vdd raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3912.71fF
C12319 BU_3VX2_51|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.71fF
C12320 BU_3VX2_50|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.70fF
C12321 BU_3VX2_49|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.28fF
C12322 BU_3VX2_48|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.92fF
C12323 BU_3VX2_47|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.94fF
C12324 adc0_data<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.88fF
C12325 BU_3VX2_46|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.34fF
C12326 BU_3VX2_45|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.66fF
C12327 BU_3VX2_44|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.39fF
C12328 BU_3VX2_43|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.46fF
C12329 BU_3VX2_42|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.25fF
C12330 LS_3VX2_20|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.65fF
C12331 LS_3VX2_21|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.90fF
C12332 LS_3VX2_27|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.70fF
C12333 BU_3VX2_52|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.92fF
C12334 BU_3VX2_53|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.82fF
C12335 BU_3VX2_54|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.10fF
C12336 BU_3VX2_55|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.13fF
C12337 BU_3VX2_56|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.16fF
C12338 BU_3VX2_57|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.26fF
C12339 BU_3VX2_58|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.89fF
C12340 BU_3VX2_59|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.08fF
C12341 BU_3VX2_60|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.77fF
C12342 BU_3VX2_61|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.02fF
C12343 BU_3VX2_62|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.10fF
C12344 LS_3VX2_15|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.98fF
C12345 LS_3VX2_16|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.73fF
C12346 LS_3VX2_17|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.74fF
C12347 AMUX4_3V_0|SEL[1] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.29fF
C12348 AMUX4_3V_0|SEL[0] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -9.06fF
C12349 AMUX4_3V_4|AIN2 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 10.68fF
C12350 BU_3VX2_42|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.04fF
C12351 LS_3VX2_27|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.03fF
C12352 LS_3VX2_21|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.01fF
C12353 LS_3VX2_20|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.08fF
C12354 BU_3VX2_43|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.34fF
C12355 BU_3VX2_44|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.60fF
C12356 BU_3VX2_45|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.87fF
C12357 BU_3VX2_46|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.39fF
C12358 BU_3VX2_41|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.39fF
C12359 BU_3VX2_47|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.48fF
C12360 BU_3VX2_48|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.49fF
C12361 BU_3VX2_49|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.51fF
C12362 BU_3VX2_50|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.44fF
C12363 BU_3VX2_51|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.44fF
C12364 AMUX4_3V_0|AOUT raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.91fF
C12365 AMUX4_3V_1|SEL[1] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -11.75fF
C12366 AMUX4_3V_1|SEL[0] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -9.74fF
C12367 comp_inp raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 54.70fF
C12368 AMUX4_3V_4|AIN3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 10.18fF
C12369 BU_3VX2_62|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.04fF
C12370 LS_3VX2_17|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.90fF
C12371 LS_3VX2_16|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.95fF
C12372 LS_3VX2_15|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.00fF
C12373 BU_3VX2_61|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.44fF
C12374 BU_3VX2_60|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12375 BU_3VX2_59|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12376 BU_3VX2_58|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12377 BU_3VX2_57|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12378 BU_3VX2_56|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12379 BU_3VX2_55|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12380 BU_3VX2_54|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.37fF
C12381 BU_3VX2_53|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.49fF
C12382 BU_3VX2_52|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.53fF
C12383 VDD3V3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 584.44fF
C12384 AMUX4_3V_1|AOUT raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.54fF
C12385 BU_3VX2_17|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.16fF
C12386 BU_3VX2_8|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.62fF
C12387 BU_3VX2_20|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.42fF
C12388 BU_3VX2_10|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.18fF
C12389 BU_3VX2_67|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.15fF
C12390 BU_3VX2_22|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.86fF
C12391 BU_3VX2_9|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.01fF
C12392 BU_3VX2_7|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -6.72fF
C12393 BU_3VX2_18|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.86fF
C12394 BU_3VX2_30|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.11fF
C12395 BU_3VX2_33|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.28fF
C12396 BU_3VX2_69|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.40fF
C12397 BU_3VX2_65|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.39fF
C12398 BU_3VX2_31|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.68fF
C12399 BU_3VX2_5|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.50fF
C12400 BU_3VX2_64|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.60fF
C12401 BU_3VX2_68|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.27fF
C12402 AMUX4_3V_4|SEL[1] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.74fF
C12403 AMUX4_3V_3|SEL[0] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.81fF
C12404 BU_3VX2_36|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.82fF
C12405 AMUX4_3V_4|SEL[0] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.91fF
C12406 BU_3VX2_4|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.60fF
C12407 LS_3VX2_23|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.19fF
C12408 BU_3VX2_11|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.58fF
C12409 BU_3VX2_32|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.58fF
C12410 BU_3VX2_70|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.15fF
C12411 BU_3VX2_3|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.50fF
C12412 BU_3VX2_37|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.45fF
C12413 BU_3VX2_14|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.41fF
C12414 raven_soc_0|ram_rdata<16> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.33fF
C12415 raven_soc_0|ram_rdata<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.80fF
C12416 raven_soc_0|ram_addr<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.01fF
C12417 raven_soc_0|ram_rdata<17> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.42fF
C12418 raven_soc_0|ram_rdata<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.48fF
C12419 raven_soc_0|ram_rdata<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.11fF
C12420 raven_soc_0|ram_wdata<31> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.26fF
C12421 raven_soc_0|ram_wdata<27> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.39fF
C12422 raven_soc_0|ram_wdata<29> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.28fF
C12423 raven_soc_0|ram_wdata<22> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.99fF
C12424 raven_soc_0|ram_wdata<25> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.42fF
C12425 raven_soc_0|ram_wdata<21> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.28fF
C12426 raven_soc_0|ram_wdata<19> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.19fF
C12427 raven_soc_0|ram_wdata<26> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.78fF
C12428 raven_soc_0|ram_wdata<17> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.78fF
C12429 raven_soc_0|ram_rdata<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.85fF
C12430 raven_soc_0|ram_wdata<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.79fF
C12431 raven_soc_0|ram_wdata<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.02fF
C12432 raven_soc_0|ram_wdata<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.31fF
C12433 raven_soc_0|ram_rdata<25> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.49fF
C12434 raven_soc_0|ram_wdata<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.13fF
C12435 raven_soc_0|ram_wdata<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.06fF
C12436 raven_soc_0|irq_pin raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.64fF
C12437 raven_soc_0|ram_rdata<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.07fF
C12438 raven_soc_0|ram_wdata<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.04fF
C12439 raven_soc_0|ram_wdata<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.05fF
C12440 raven_soc_0|ram_rdata<23> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.10fF
C12441 raven_soc_0|ram_rdata<19> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.17fF
C12442 raven_soc_0|ram_rdata<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.50fF
C12443 raven_soc_0|ram_rdata<20> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.00fF
C12444 raven_soc_0|ram_rdata<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.29fF
C12445 raven_soc_0|ram_rdata<28> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.71fF
C12446 raven_soc_0|flash_clk raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.27fF
C12447 raven_soc_0|flash_io1_oeb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.09fF
C12448 raven_soc_0|flash_io0_do raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.45fF
C12449 raven_soc_0|flash_io2_di raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.77fF
C12450 raven_soc_0|flash_io0_di raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.90fF
C12451 raven_soc_0|flash_io3_di raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.97fF
C12452 raven_soc_0|flash_io0_oeb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.47fF
C12453 raven_soc_0|flash_io3_oeb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.66fF
C12454 raven_soc_0|flash_io1_di raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.25fF
C12455 raven_soc_0|flash_io2_oeb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.63fF
C12456 raven_soc_0|flash_io1_do raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.08fF
C12457 raven_soc_0|flash_io2_do raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.78fF
C12458 raven_soc_0|flash_io3_do raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.65fF
C12459 raven_soc_0|gpio_out<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 26.61fF
C12460 raven_soc_0|gpio_in<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.96fF
C12461 raven_soc_0|gpio_in<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 16.97fF
C12462 raven_soc_0|gpio_in<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.22fF
C12463 raven_soc_0|gpio_in<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.63fF
C12464 raven_soc_0|gpio_in<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.47fF
C12465 raven_soc_0|gpio_in<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.65fF
C12466 raven_soc_0|gpio_in<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.82fF
C12467 raven_soc_0|gpio_in<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.15fF
C12468 raven_soc_0|gpio_in<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.90fF
C12469 raven_soc_0|gpio_in<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 12.22fF
C12470 raven_soc_0|gpio_pullup<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.71fF
C12471 raven_soc_0|ext_clk raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.02fF
C12472 BU_3VX2_40|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -10.77fF
C12473 raven_soc_0|ram_rdata<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.36fF
C12474 raven_soc_0|ram_rdata<31> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -6.68fF
C12475 raven_soc_0|ram_wdata<24> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.75fF
C12476 raven_soc_0|ram_wdata<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.09fF
C12477 raven_soc_0|ram_wdata<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.39fF
C12478 raven_soc_0|ram_rdata<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.58fF
C12479 raven_soc_0|ram_rdata<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.06fF
C12480 raven_soc_0|ram_addr<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -8.80fF
C12481 raven_soc_0|ram_wdata<20> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.83fF
C12482 raven_soc_0|ram_addr<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.07fF
C12483 raven_soc_0|ram_addr<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.18fF
C12484 raven_soc_0|ram_rdata<30> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 9.50fF
C12485 raven_soc_0|ram_rdata<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.73fF
C12486 raven_soc_0|ram_wdata<23> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.87fF
C12487 raven_soc_0|ram_rdata<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.28fF
C12488 raven_soc_0|ram_rdata<24> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.59fF
C12489 raven_soc_0|ram_rdata<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.75fF
C12490 raven_soc_0|ram_rdata<18> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.18fF
C12491 raven_soc_0|ram_rdata<21> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.07fF
C12492 raven_soc_0|ram_rdata<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.09fF
C12493 raven_soc_0|ram_wdata<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.92fF
C12494 raven_soc_0|ram_rdata<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.48fF
C12495 raven_soc_0|ram_rdata<22> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.40fF
C12496 LS_3VX2_18|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.73fF
C12497 raven_soc_0|ser_tx raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.84fF
C12498 LS_3VX2_2|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.49fF
C12499 BU_3VX2_1|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.15fF
C12500 LS_3VX2_19|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -8.33fF
C12501 LS_3VX2_22|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.93fF
C12502 BU_3VX2_21|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.85fF
C12503 BU_3VX2_66|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.61fF
C12504 BU_3VX2_2|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.31fF
C12505 BU_3VX2_13|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.39fF
C12506 BU_3VX2_38|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.67fF
C12507 BU_3VX2_12|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.26fF
C12508 BU_3VX2_15|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.10fF
C12509 BU_3VX2_6|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.07fF
C12510 BU_3VX2_19|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.62fF
C12511 BU_3VX2_16|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.08fF
C12512 BU_3VX2_73|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.83fF
C12513 BU_3VX2_35|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.79fF
C12514 BU_3VX2_71|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -14.70fF
C12515 raven_soc_0|gpio_outenb<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.29fF
C12516 raven_soc_0|gpio_out<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.08fF
C12517 raven_soc_0|gpio_in<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.15fF
C12518 raven_soc_0|gpio_outenb<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.44fF
C12519 raven_soc_0|gpio_pullup<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 14.53fF
C12520 raven_soc_0|gpio_outenb<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.86fF
C12521 raven_soc_0|gpio_out<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.23fF
C12522 raven_soc_0|gpio_out<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.64fF
C12523 raven_soc_0|gpio_pullup<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.63fF
C12524 raven_soc_0|gpio_pullup<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.38fF
C12525 raven_soc_0|gpio_pulldown<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.36fF
C12526 raven_soc_0|gpio_pulldown<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.58fF
C12527 raven_soc_0|gpio_pulldown<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.03fF
C12528 AMUX4_3V_3|SEL[1] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.69fF
C12529 raven_soc_0|ram_addr<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.34fF
C12530 raven_soc_0|ram_addr<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.03fF
C12531 raven_soc_0|ram_addr<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.36fF
C12532 raven_soc_0|ram_addr<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.69fF
C12533 raven_soc_0|ram_addr<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.83fF
C12534 raven_soc_0|ram_addr<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.98fF
C12535 raven_soc_0|ram_rdata<29> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 9.24fF
C12536 raven_soc_0|ram_rdata<27> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.17fF
C12537 raven_soc_0|ram_rdata<26> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.66fF
C12538 raven_soc_0|ram_rdata<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.00fF
C12539 raven_soc_0|ram_wdata<30> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.96fF
C12540 raven_soc_0|ram_wdata<28> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.71fF
C12541 raven_soc_0|ram_wdata<18> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.54fF
C12542 raven_soc_0|ram_wdata<16> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.66fF
C12543 raven_soc_0|ram_wdata<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.21fF
C12544 raven_soc_0|ram_wdata<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.10fF
C12545 raven_soc_0|ram_wdata<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.25fF
C12546 raven_soc_0|ram_wdata<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.13fF
C12547 raven_soc_0|ram_wdata<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.76fF
C12548 raven_soc_0|ram_wdata<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.19fF
C12549 raven_soc_0|ram_wenb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.38fF
C12550 raven_soc_0|flash_csb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -22.67fF
C12551 raven_soc_0|gpio_out<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.61fF
C12552 raven_soc_0|gpio_out<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -9.08fF
C12553 raven_soc_0|gpio_out<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.46fF
C12554 raven_soc_0|gpio_out<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.38fF
C12555 raven_soc_0|gpio_out<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.81fF
C12556 raven_soc_0|gpio_out<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.02fF
C12557 raven_soc_0|gpio_out<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.21fF
C12558 raven_soc_0|gpio_outenb<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 28.97fF
C12559 raven_soc_0|gpio_outenb<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -6.51fF
C12560 raven_soc_0|gpio_outenb<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.60fF
C12561 raven_soc_0|gpio_outenb<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.03fF
C12562 raven_soc_0|gpio_outenb<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.75fF
C12563 raven_soc_0|gpio_outenb<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.89fF
C12564 raven_soc_0|gpio_outenb<6> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.43fF
C12565 raven_soc_0|gpio_outenb<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.58fF
C12566 raven_soc_0|gpio_pullup<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 49.17fF
C12567 raven_soc_0|gpio_pullup<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.75fF
C12568 raven_soc_0|gpio_pullup<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.40fF
C12569 raven_soc_0|gpio_pullup<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -8.82fF
C12570 raven_soc_0|gpio_pullup<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.49fF
C12571 raven_soc_0|gpio_pullup<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.64fF
C12572 raven_soc_0|gpio_pullup<7> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.10fF
C12573 raven_soc_0|gpio_pullup<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.02fF
C12574 raven_soc_0|gpio_pullup<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.20fF
C12575 raven_soc_0|gpio_pulldown<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.47fF
C12576 raven_soc_0|gpio_pulldown<5> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.70fF
C12577 raven_soc_0|gpio_pulldown<8> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.65fF
C12578 raven_soc_0|gpio_pulldown<9> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.53fF
C12579 raven_soc_0|gpio_pulldown<10> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -7.33fF
C12580 raven_soc_0|gpio_pulldown<11> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.89fF
C12581 raven_soc_0|gpio_pulldown<12> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.11fF
C12582 raven_soc_0|gpio_pulldown<13> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.68fF
C12583 raven_soc_0|gpio_pulldown<14> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 13.84fF
C12584 raven_soc_0|gpio_pulldown<15> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.45fF
C12585 raven_soc_0|ser_rx raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 4.14fF
C12586 BU_3VX2_0|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -27.45fF
C12587 BU_3VX2_63|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -11.51fF
C12588 AMUX2_3V_0|SEL raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.57fF
C12589 LS_3VX2_3|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -15.25fF
C12590 LS_3VX2_13|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.34fF
C12591 LS_3VX2_12|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.68fF
C12592 LS_3VX2_11|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.70fF
C12593 LS_3VX2_10|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.20fF
C12594 LS_3VX2_9|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -9.96fF
C12595 LS_3VX2_14|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -7.12fF
C12596 LS_3VX2_8|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.69fF
C12597 LS_3VX2_7|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.77fF
C12598 LS_3VX2_6|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.67fF
C12599 LS_3VX2_5|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.00fF
C12600 LS_3VX2_4|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -9.04fF
C12601 LS_3VX2_24|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.50fF
C12602 LS_3VX2_24|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -10.20fF
C12603 LS_3VX2_14|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.90fF
C12604 LS_3VX2_4|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.39fF
C12605 LS_3VX2_9|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.62fF
C12606 LS_3VX2_5|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.58fF
C12607 LS_3VX2_10|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.40fF
C12608 LS_3VX2_6|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.33fF
C12609 LS_3VX2_11|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.53fF
C12610 LS_3VX2_7|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.60fF
C12611 LS_3VX2_12|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.74fF
C12612 LS_3VX2_8|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.72fF
C12613 LS_3VX2_13|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.41fF
C12614 AMUX2_3V_0|AOUT raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.71fF
C12615 acsoc02_3v3_0|CS_8U raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.04fF
C12616 acsoc02_3v3_0|CS_4U raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.04fF
C12617 LS_3VX2_19|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.76fF
C12618 aopac01_3v3_0|IB raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.14fF
C12619 LS_3VX2_22|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.31fF
C12620 BU_3VX2_73|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.90fF
C12621 BU_3VX2_40|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.12fF
C12622 BU_3VX2_35|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.92fF
C12623 BU_3VX2_38|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.66fF
C12624 BU_3VX2_37|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.17fF
C12625 BU_3VX2_2|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.86fF
C12626 BU_3VX2_11|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -7.47fF
C12627 BU_3VX2_12|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.14fF
C12628 BU_3VX2_13|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.41fF
C12629 BU_3VX2_14|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.39fF
C12630 BU_3VX2_15|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.78fF
C12631 BU_3VX2_16|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.56fF
C12632 BU_3VX2_17|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.59fF
C12633 BU_3VX2_18|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.43fF
C12634 BU_3VX2_19|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.35fF
C12635 BU_3VX2_20|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.42fF
C12636 BU_3VX2_21|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.21fF
C12637 BU_3VX2_22|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.24fF
C12638 BU_3VX2_23|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.35fF
C12639 BU_3VX2_24|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.22fF
C12640 BU_3VX2_25|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.82fF
C12641 BU_3VX2_26|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.83fF
C12642 BU_3VX2_27|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.28fF
C12643 BU_3VX2_28|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.22fF
C12644 BU_3VX2_29|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.14fF
C12645 BU_3VX2_33|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 5.83fF
C12646 BU_3VX2_36|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.78fF
C12647 BU_3VX2_64|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.07fF
C12648 BU_3VX2_65|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.74fF
C12649 BU_3VX2_66|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.11fF
C12650 BU_3VX2_67|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.75fF
C12651 BU_3VX2_68|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.16fF
C12652 BU_3VX2_69|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.48fF
C12653 BU_3VX2_70|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.57fF
C12654 BU_3VX2_6|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.06fF
C12655 raven_spi_0|SDI raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.70fF
C12656 BU_3VX2_10|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.14fF
C12657 raven_spi_0|SDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.04fF
C12658 raven_spi_0|CSB raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.68fF
C12659 BU_3VX2_63|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.19fF
C12660 BU_3VX2_71|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.01fF
C12661 LS_3VX2_3|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.06fF
C12662 BU_3VX2_4|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.44fF
C12663 BU_3VX2_5|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.63fF
C12664 BU_3VX2_9|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.54fF
C12665 BU_3VX2_8|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.58fF
C12666 BU_3VX2_7|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -1.30fF
C12667 BU_3VX2_3|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.06fF
C12668 aporc02_3v3_0|PORB raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.07fF
C12669 BU_3VX2_0|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.65fF
C12670 BU_3VX2_1|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.55fF
C12671 LS_3VX2_2|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.04fF
C12672 acsoc01_3v3_0|CS3_200N raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.05fF
C12673 acsoc01_3v3_0|CS2_200N raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.05fF
C12674 BU_3VX2_32|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 17.74fF
C12675 LS_3VX2_23|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.84fF
C12676 acmpc01_3v3_0|IBN raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.84fF
C12677 LS_3VX2_18|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.33fF
C12678 XSPRAM_1024X32_M8P_0|RDY raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12679 AMUX4_3V_4|AOUT raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 7.57fF
C12680 AMUX4_3V_3|AOUT raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.38fF
C12681 LOGIC1_3V_0|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.24fF
C12682 LOGIC1_3V_1|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.24fF
C12683 LOGIC1_3V_2|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.24fF
C12684 LOGIC1_3V_3|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.24fF
C12685 LOGIC0_3V_0|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.11fF
C12686 LOGIC0_3V_1|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.10fF
C12687 LOGIC0_3V_2|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.04fF
C12688 LOGIC0_3V_3|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.25fF
C12689 XI raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.82fF
C12690 XO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -3.85fF
C12691 SDO raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.65fF
C12692 SCK raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 37.87fF
C12693 CSB raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 12.42fF
C12694 SDI raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 18.78fF
C12695 gpio[15] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 33.10fF
C12696 ser_rx raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 8.32fF
C12697 ser_tx raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 36.03fF
C12698 irq raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 43.71fF
C12699 gpio[14] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 42.34fF
C12700 gpio[13] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.55fF
C12701 comp_inn raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 45.54fF
C12702 gpio[12] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.55fF
C12703 gpio[11] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.06fF
C12704 VSS raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 45.90fF
C12705 gpio[10] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 31.51fF
C12706 gpio[9] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.45fF
C12707 gpio[8] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.07fF
C12708 gpio[7] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 41.95fF
C12709 gpio[6] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 41.76fF
C12710 gpio[5] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 39.67fF
C12711 gpio[4] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 25.15fF
C12712 gpio[3] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 41.02fF
C12713 adc1_in raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 41.83fF
C12714 adc0_in raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.97fF
C12715 gpio[0] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 6.15fF
C12716 gpio[1] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -4.82fF
C12717 gpio[2] raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -66.11fF
C12718 IN_3VX2_1|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.02fF
C12719 raven_soc_0|gpio_pullup<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -8.48fF
C12720 AMUX4_3V_0|AIN1 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 15.12fF
C12721 raven_soc_0|gpio_out<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.83fF
C12722 AMUX4_3V_1|AIN1 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -2.56fF
C12723 raven_soc_0|gpio_out<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.36fF
C12724 raven_soc_0|gpio_in<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.14fF
C12725 raven_soc_0|gpio_out<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.89fF
C12726 raven_soc_0|gpio_in<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -7.41fF
C12727 raven_soc_0|gpio_in<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.16fF
C12728 flash_io2 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 42.17fF
C12729 flash_clk raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 10.83fF
C12730 raven_soc_0|gpio_pulldown<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.57fF
C12731 raven_soc_0|gpio_outenb<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.03fF
C12732 flash_io1 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 40.44fF
C12733 raven_soc_0|gpio_pullup<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.47fF
C12734 flash_io0 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 43.32fF
C12735 raven_soc_0|gpio_outenb<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.43fF
C12736 raven_soc_0|gpio_out<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.76fF
C12737 raven_soc_0|gpio_pulldown<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.34fF
C12738 adc_high raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 11.81fF
C12739 flash_io3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 42.65fF
C12740 raven_soc_0|gpio_in<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -12.87fF
C12741 raven_spi_0|sdo_enb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.09fF
C12742 raven_soc_0|gpio_in<2> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.92fF
C12743 raven_soc_0|gpio_outenb<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 1.29fF
C12744 XCLK raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 36.28fF
C12745 raven_soc_0|gpio_out<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.24fF
C12746 raven_soc_0|gpio_outenb<4> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.91fF
C12747 adc_low raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 51.25fF
C12748 raven_soc_0|gpio_outenb<3> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -0.75fF
C12749 raven_soc_0|gpio_pulldown<1> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -5.67fF
C12750 BU_3VX2_31|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -20.62fF
C12751 flash_csb raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 41.59fF
C12752 analog_out raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 18.10fF
C12753 AMUX4_3V_4|AIN1 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.71fF
C12754 raven_soc_0|gpio_pullup<0> raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 2.15fF
C12755 IN_3VX2_1|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# -35.09fF
C12756 LOGIC0_3V_4|Q raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 689.31fF
C12757 BU_3VX2_72|A raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.71fF
C12758 raven_padframe_0|BBCUD4F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12759 raven_padframe_0|BBCUD4F_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12760 raven_padframe_0|FILLER02F_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12761 raven_padframe_0|FILLER20F_3|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12762 raven_padframe_0|GNDORPADF_7|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.83fF
C12763 raven_padframe_0|FILLER10F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12764 raven_padframe_0|FILLER02F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12765 raven_padframe_0|FILLER20F_5|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12766 raven_padframe_0|BBCUD4F_3|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12767 raven_padframe_0|BBCUD4F_4|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12768 raven_padframe_0|BBCUD4F_6|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12769 raven_padframe_0|BBCUD4F_5|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12770 raven_padframe_0|BBCUD4F_7|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12771 raven_padframe_0|BBCUD4F_8|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12772 raven_padframe_0|BBCUD4F_9|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12773 raven_padframe_0|BBCUD4F_10|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12774 raven_padframe_0|BBCUD4F_11|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12775 raven_padframe_0|BBCUD4F_13|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12776 raven_padframe_0|BBCUD4F_12|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12777 raven_padframe_0|BBCUD4F_14|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.03fF
C12778 raven_padframe_0|GNDORPADF_3|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.81fF
C12779 raven_padframe_0|ICF_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12780 raven_padframe_0|BT4F_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12781 raven_padframe_0|BT4F_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12782 raven_padframe_0|BBC4F_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12783 raven_padframe_0|BBC4F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12784 raven_padframe_0|BBC4F_3|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12785 raven_padframe_0|BBC4F_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12786 raven_padframe_0|FILLER40F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12787 raven_padframe_0|POWERCUTVDD3FC_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12788 raven_padframe_0|VDDPADFC_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12789 raven_padframe_0|BT4FC_0|VDD3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.05fF
C12790 raven_padframe_0|BT4FC_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12791 raven_padframe_0|ICFC_2|VDD3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.05fF
C12792 raven_padframe_0|ICFC_2|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12793 raven_padframe_0|ICFC_1|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12794 raven_padframe_0|ICFC_1|VDD3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.05fF
C12795 raven_padframe_0|ICFC_0|VDD3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.08fF
C12796 raven_padframe_0|ICFC_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12797 raven_padframe_0|FILLER20FC_0|VDD3 raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.05fF
C12798 raven_padframe_0|FILLER20FC_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12799 raven_padframe_0|FILLER20F_8|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12800 raven_padframe_0|POWERCUTVDD3FC_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12801 raven_padframe_0|BBCUD4F_15|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12802 raven_padframe_0|GNDORPADF_5|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
C12803 VDD raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 3.08fF
C12804 raven_padframe_0|FILLER20F_0|VDDR raven_padframe_0|CORNERESDF_1|w_n1073741817_n1073741817# 0.02fF
.ends

