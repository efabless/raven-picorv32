module acsoc01_3v3 ( CS1_200N, CS0_200N, EN, VDDA, VSSA, CS2_200N, CS3_200N
);

  input EN;
  input VSSA;
  input VDDA;
  input CS1_200N;
  input CS3_200N;
  input CS2_200N;
  input CS0_200N;

  wire real CS1_200N;
  wire real CS3_200N;
  wire real CS2_200N;
  wire real CS0_200N;

endmodule
