module analog_isource2_3v3 ( CS_2U, CS_1U, EN, VDDA, VSSA, CS_4U, CS_8U );

  input EN;
  input VSSA;
  input VDDA;
  input CS_4U;
  input CS_1U;
  input CS_8U;
  input CS_2U;

  wire real VSSA, VDDA;
  wire real CS_4U;
  wire real CS_1U;
  wire real CS_8U;
  wire real CS_2U;

  

endmodule
