* NGSPICE file created from raven.ext - technology: EFXH018D

* Black-box entry subcircuit for CORNERESDF abstract view
.subckt CORNERESDF GNDR VDDR VDD VDDO GNDO
.ends

* Black-box entry subcircuit for FILLER01F abstract view
.subckt FILLER01F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for FILLER10F abstract view
.subckt FILLER10F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for FILLER20F abstract view
.subckt FILLER20F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for FILLER50F abstract view
.subckt FILLER50F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for VDDPADF abstract view
.subckt VDDPADF VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for VDDORPADF abstract view
.subckt VDDORPADF VDDOR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for GNDORPADF abstract view
.subckt GNDORPADF VDDO VDDR VDD GNDOR
.ends

* Black-box entry subcircuit for ICF abstract view
.subckt ICF PO PI Y PAD VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for BT4F abstract view
.subckt BT4F EN A PAD VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for BBC4F abstract view
.subckt BBC4F EN A Y PO PI PAD VDDO GNDO GNDR VDDR VDD
.ends

* Black-box entry subcircuit for FILLER40F abstract view
.subckt FILLER40F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for POWERCUTVDD3FC abstract view
.subckt POWERCUTVDD3FC VDDO VDDR GNDR GNDO
.ends

* Black-box entry subcircuit for VDDPADFC abstract view
.subckt VDDPADFC VDDO VDDR GNDR GNDO VDD3
.ends

* Black-box entry subcircuit for BT4FC abstract view
.subckt BT4FC EN A PAD VDDO VDDR GNDR GNDO VDD3
.ends

* Black-box entry subcircuit for ICFC abstract view
.subckt ICFC PO PI Y PAD VDDO VDDR GNDR GNDO VDD3
.ends

* Black-box entry subcircuit for FILLER20FC abstract view
.subckt FILLER20FC VDDO VDDR GNDR GNDO VDD3
.ends

* Black-box entry subcircuit for BBCUD4F abstract view
.subckt BBCUD4F EN A Y PO PI PUEN PDEN PAD VDDO GNDO GNDR VDDR VDD
.ends

* Black-box entry subcircuit for APR00DF abstract view
.subckt APR00DF PAD VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for aregc01_3v3 abstract view
.subckt aregc01_3v3 OUT EN VIN3 ENB VDD VDDR GNDR GNDO VDDO
.ends

* Black-box entry subcircuit for FILLER02F abstract view
.subckt FILLER02F VDDO VDDR GNDR GNDO VDD
.ends

* Black-box entry subcircuit for axtoc02_3v3 abstract view
.subckt axtoc02_3v3 GNDO VDDO GNDR VDDR VDD XI XO CLK EN
.ends

.subckt raven_padframe BBCUD4F_0/PI BBCUD4F_4/EN gpio<10> VDD3V3 XCLK comp_inn BBCUD4F_8/PDEN
+ VSS BBCUD4F_5/Y BBCUD4F_9/PUEN BBCUD4F_2/A ICF_2/PI comp_inp SCK gpio<9> BBC4F_3/A
+ BBCUD4F_14/PI BBCUD4F_0/EN flash_io0 comp_inp BBCUD4F_7/PI BBC4F_1/PI BBCUD4F_0/PDEN
+ ICF_1/Y gpio<14> BBCUD4F_13/Y BBCUD4F_1/PUEN BT4F_2/A BBCUD4F_13/PDEN BBCUD4F_10/A
+ VDD1V8 gpio<2> BBCUD4F_14/PUEN BBCUD4F_9/Y VDD3V3 BT4F_2/EN BBCUD4F_6/A irq BBCUD4F_10/PI
+ BBCUD4F_7/PDEN BBCUD4F_8/PUEN BBCUD4F_0/Y BBCUD4F_14/EN BBCUD4F_3/PI BBC4F_1/EN
+ BBCUD4F_7/EN BBC4F_1/Y ICFC_0/PI APR00DF_3/PAD BBCUD4F_14/A BT4FC_0/A gpio<6> BT4FC_0/EN
+ BBCUD4F_12/PDEN BBCUD4F_0/PUEN VSS BBCUD4F_13/PUEN axtoc02_3v3_0/CLK BBCUD4F_10/EN
+ BBCUD4F_4/Y BBCUD4F_3/EN VSS gpio<11> BBCUD4F_1/A SDI BBC4F_2/A BBCUD4F_6/PDEN BBCUD4F_7/PUEN
+ VDD3V3 ICF_1/PI XCLK ICF_0/Y BBCUD4F_12/Y adc0_in BT4F_1/A ICFC_0/VDD3 BBCUD4F_13/PI
+ BBCUD4F_8/Y axtoc02_3v3_0/EN w_n1073741817_n1073741817# BBCUD4F_6/PI BBC4F_0/PI
+ BBCUD4F_5/A flash_io1 BBCUD4F_11/PDEN BBCUD4F_12/PUEN gpio<15> gpio<3> BBC4F_0/Y
+ BT4F_1/EN aregc01_3v3_1/EN BBCUD4F_5/PDEN BBCUD4F_6/PUEN ICFC_2/Y BBCUD4F_13/A BBCUD4F_13/EN
+ BBCUD4F_2/PI SDO BBC4F_0/EN BBCUD4F_6/EN BBCUD4F_9/A ser_tx APR00DF_4/PAD BBCUD4F_3/Y
+ aregc01_3v3_0/ENB gpio<7> BBCUD4F_0/A BBCUD4F_10/PDEN adc1_in BBC4F_1/A BBCUD4F_11/PUEN
+ BBCUD4F_2/EN BBCUD4F_9/PI BBC4F_3/PI gpio<12> BBCUD4F_11/Y gpio<0> BT4F_0/A BBCUD4F_5/PUEN
+ BBCUD4F_4/PDEN BBCUD4F_7/Y flash_csb BBCUD4F_4/A ICF_0/PI VSS BBCUD4F_12/PI adc1_in
+ BBCUD4F_5/PI VDD3V3 ICFC_2/PI BBC4F_3/EN BBCUD4F_9/EN BBCUD4F_10/PUEN flash_io3
+ BBCUD4F_15/Y VDD3V3 aregc01_3v3_0/OUT BBCUD4F_12/A ICFC_1/Y gpio<4> BT4F_0/EN aregc01_3v3_0/EN
+ BBCUD4F_8/A flash_clk BBCUD4F_3/PDEN BBCUD4F_4/PUEN BBCUD4F_12/EN BBCUD4F_2/Y BBCUD4F_1/PI
+ BBC4F_3/Y flash_io0 VDD1V8 BBCUD4F_5/EN BBC4F_0/A flash_io1 comp_inn XI adc0_in
+ flash_io2 gpio<8> aregc01_3v3_1/ENB BBCUD4F_10/Y flash_io3 BBCUD4F_6/Y BBCUD4F_15/PI
+ BBCUD4F_1/EN BBCUD4F_8/PI BBC4F_2/PI BBCUD4F_3/A gpio<13> VDD1V8 BBCUD4F_3/PUEN
+ BBCUD4F_2/PDEN gpio<1> BBCUD4F_15/PDEN aregc01_3v3_1/VIN3 CSB ICF_2/Y BBCUD4F_14/Y
+ BBCUD4F_11/PI ICFC_0/Y flash_clk BBCUD4F_11/A BBCUD4F_9/PDEN BBCUD4F_15/EN VSS BBCUD4F_4/PI
+ ser_rx BBCUD4F_8/EN BBC4F_2/EN ICFC_1/PI APR00DF_2/PAD BBCUD4F_7/A XO flash_io2
+ gpio<5> BBCUD4F_1/Y VSS aregc01_3v3_1/OUT BBC4F_2/Y BBCUD4F_1/PDEN VDD3V3 BBCUD4F_14/PDEN
+ BBCUD4F_15/PUEN flash_csb BBCUD4F_2/PUEN aregc01_3v3_0/VIN3 BBCUD4F_11/EN BBCUD4F_15/A
XCORNERESDF_3 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER01F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER01F
XFILLER10F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER10F
XFILLER20F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XFILLER50F_2 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XVDDPADF_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 VDDPADF
XVDDORPADF_4 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_3 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XICF_2 ICF_2/PO ICF_2/PI ICF_2/Y XCLK VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XBT4F_1 BT4F_1/EN BT4F_1/A flash_clk VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XBT4F_2 BT4F_2/EN BT4F_2/A flash_csb VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XBBC4F_0 BBC4F_0/EN BBC4F_0/A BBC4F_0/Y BBC4F_0/PO BBC4F_0/PI flash_io0 VDD3V3 VSS
+ VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_1 BBC4F_1/EN BBC4F_1/A BBC4F_1/Y BBC4F_1/PO BBC4F_1/PI flash_io1 VDD3V3 VSS
+ VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_3 BBC4F_3/EN BBC4F_3/A BBC4F_3/Y BBC4F_3/PO BBC4F_3/PI flash_io2 VDD3V3 VSS
+ VSS VDD3V3 VDD1V8 BBC4F
XBBC4F_2 BBC4F_2/EN BBC4F_2/A BBC4F_2/Y BBC4F_2/PO BBC4F_2/PI flash_io3 VDD3V3 VSS
+ VSS VDD3V3 VDD1V8 BBC4F
XFILLER40F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER40F
XPOWERCUTVDD3FC_1 VDD3V3 VDD3V3 VSS VSS POWERCUTVDD3FC
XVDDPADFC_0 VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 VDDPADFC
XBT4FC_0 BT4FC_0/EN BT4FC_0/A SDO VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 BT4FC
XICFC_2 ICFC_2/PO ICFC_2/PI ICFC_2/Y SCK VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 ICFC
XICFC_1 ICFC_1/PO ICFC_1/PI ICFC_1/Y CSB VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 ICFC
XFILLER20FC_0 VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 FILLER20FC
XICFC_0 ICFC_0/PO ICFC_0/PI ICFC_0/Y SDI VDD3V3 VDD3V3 VSS VSS ICFC_0/VDD3 ICFC
XPOWERCUTVDD3FC_0 VDD3V3 VDD3V3 VSS VSS POWERCUTVDD3FC
XFILLER20F_8 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XBBCUD4F_15 BBCUD4F_15/EN BBCUD4F_15/A BBCUD4F_15/Y BBCUD4F_15/PO BBCUD4F_15/PI BBCUD4F_15/PUEN
+ BBCUD4F_15/PDEN gpio<15> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XGNDORPADF_5 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER20F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_2 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER20F_7 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XICF_0 ICF_0/PO ICF_0/PI ICF_0/Y ser_rx VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XBT4F_0 BT4F_0/EN BT4F_0/A ser_tx VDD3V3 VDD3V3 VSS VSS VDD1V8 BT4F
XICF_1 ICF_1/PO ICF_1/PI ICF_1/Y irq VDD3V3 VDD3V3 VSS VSS VDD1V8 ICF
XAPR00DF_6 comp_inp VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_5 comp_inn VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XFILLER50F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XGNDORPADF_0 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XVDDORPADF_0 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XVDDPADF_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 VDDPADF
XFILLER20F_6 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XGNDORPADF_2 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER50F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER50F
XGNDORPADF_6 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XVDDORPADF_2 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XFILLER01F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER01F
XBBCUD4F_14 BBCUD4F_14/EN BBCUD4F_14/A BBCUD4F_14/Y BBCUD4F_14/PO BBCUD4F_14/PI BBCUD4F_14/PUEN
+ BBCUD4F_14/PDEN gpio<14> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_13 BBCUD4F_13/EN BBCUD4F_13/A BBCUD4F_13/Y BBCUD4F_13/PO BBCUD4F_13/PI BBCUD4F_13/PUEN
+ BBCUD4F_13/PDEN gpio<13> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_12 BBCUD4F_12/EN BBCUD4F_12/A BBCUD4F_12/Y BBCUD4F_12/PO BBCUD4F_12/PI BBCUD4F_12/PUEN
+ BBCUD4F_12/PDEN gpio<12> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_11 BBCUD4F_11/EN BBCUD4F_11/A BBCUD4F_11/Y BBCUD4F_11/PO BBCUD4F_11/PI BBCUD4F_11/PUEN
+ BBCUD4F_11/PDEN gpio<11> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_10 BBCUD4F_10/EN BBCUD4F_10/A BBCUD4F_10/Y BBCUD4F_10/PO BBCUD4F_10/PI BBCUD4F_10/PUEN
+ BBCUD4F_10/PDEN gpio<10> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_9 BBCUD4F_9/EN BBCUD4F_9/A BBCUD4F_9/Y BBCUD4F_9/PO BBCUD4F_9/PI BBCUD4F_9/PUEN
+ BBCUD4F_9/PDEN gpio<9> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_8 BBCUD4F_8/EN BBCUD4F_8/A BBCUD4F_8/Y BBCUD4F_8/PO BBCUD4F_8/PI BBCUD4F_8/PUEN
+ BBCUD4F_8/PDEN gpio<8> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_7 BBCUD4F_7/EN BBCUD4F_7/A BBCUD4F_7/Y BBCUD4F_7/PO BBCUD4F_7/PI BBCUD4F_7/PUEN
+ BBCUD4F_7/PDEN gpio<7> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
Xaregc01_3v3_1 aregc01_3v3_1/OUT aregc01_3v3_1/EN aregc01_3v3_1/VIN3 aregc01_3v3_1/ENB
+ VDD1V8 VDD3V3 VSS VSS VDD3V3 aregc01_3v3
XBBCUD4F_6 BBCUD4F_6/EN BBCUD4F_6/A BBCUD4F_6/Y BBCUD4F_6/PO BBCUD4F_6/PI BBCUD4F_6/PUEN
+ BBCUD4F_6/PDEN gpio<6> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_5 BBCUD4F_5/EN BBCUD4F_5/A BBCUD4F_5/Y BBCUD4F_5/PO BBCUD4F_5/PI BBCUD4F_5/PUEN
+ BBCUD4F_5/PDEN gpio<5> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_4 BBCUD4F_4/EN BBCUD4F_4/A BBCUD4F_4/Y BBCUD4F_4/PO BBCUD4F_4/PI BBCUD4F_4/PUEN
+ BBCUD4F_4/PDEN gpio<4> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_3 BBCUD4F_3/EN BBCUD4F_3/A BBCUD4F_3/Y BBCUD4F_3/PO BBCUD4F_3/PI BBCUD4F_3/PUEN
+ BBCUD4F_3/PDEN gpio<3> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XFILLER20F_4 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_0 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
XFILLER20F_2 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XAPR00DF_4 APR00DF_4/PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_3 APR00DF_3/PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_2 APR00DF_2/PAD VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_1 adc1_in VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XAPR00DF_0 adc0_in VDD3V3 VDD3V3 VSS VSS VDD1V8 APR00DF
XVDDORPADF_1 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_1 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
Xaregc01_3v3_0 aregc01_3v3_0/OUT aregc01_3v3_0/EN aregc01_3v3_0/VIN3 aregc01_3v3_0/ENB
+ VDD1V8 VDD3V3 VSS VSS VDD3V3 aregc01_3v3
XFILLER20F_5 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XFILLER10F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER10F
XFILLER02F_0 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER02F
XVDDORPADF_3 VDD3V3 VSS VSS VDD1V8 VDDORPADF
XGNDORPADF_7 VDD3V3 VDD3V3 VDD1V8 VSS GNDORPADF
XFILLER02F_1 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER02F
Xaxtoc02_3v3_0 VSS VDD3V3 VSS VDD3V3 VDD1V8 axtoc02_3v3_0/XI axtoc02_3v3_0/XO axtoc02_3v3_0/CLK
+ axtoc02_3v3_0/EN axtoc02_3v3
XBBCUD4F_1 BBCUD4F_1/EN BBCUD4F_1/A BBCUD4F_1/Y BBCUD4F_1/PO BBCUD4F_1/PI BBCUD4F_1/PUEN
+ BBCUD4F_1/PDEN gpio<0> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_0 BBCUD4F_0/EN BBCUD4F_0/A BBCUD4F_0/Y BBCUD4F_0/PO BBCUD4F_0/PI BBCUD4F_0/PUEN
+ BBCUD4F_0/PDEN gpio<1> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XBBCUD4F_2 BBCUD4F_2/EN BBCUD4F_2/A BBCUD4F_2/Y BBCUD4F_2/PO BBCUD4F_2/PI BBCUD4F_2/PUEN
+ BBCUD4F_2/PDEN gpio<2> VDD3V3 VSS VSS VDD3V3 VDD1V8 BBCUD4F
XFILLER20F_3 VDD3V3 VDD3V3 VSS VSS VDD1V8 FILLER20F
XCORNERESDF_1 VSS VDD3V3 VDD1V8 VDD3V3 VSS CORNERESDF
.ends

* Black-box entry subcircuit for LOGIC0_3V abstract view
.subckt LOGIC0_3V Q gnd vdd3
.ends

* Black-box entry subcircuit for LOGIC1_3V abstract view
.subckt LOGIC1_3V Q gnd vdd3
.ends

.subckt cmm5t_o8rj96 m4_n38335_n4160# m4_n6625_n4160# m4_6965_n4160# m4_n24845_n4260#
+ m4_34045_n4260# m4_11495_n4160# m4_n42965_n4260# m4_29615_n4160# m4_n24745_n4160#
+ m4_n11255_n4260# m4_20455_n4260# m4_n42865_n4160# m4_n29375_n4260# m4_38575_n4260#
+ w_n1073741817_n1073741817# m4_16025_n4160# m4_2335_n4260# m4_n11155_n4160# m4_34145_n4160#
+ m4_n29275_n4160# m4_24985_n4260# m4_n15785_n4260# m4_n33905_n4260# m4_n2195_n4260#
+ m4_20555_n4160# m4_6865_n4260# m4_n15685_n4160# m4_38675_n4160# m4_11395_n4260#
+ m4_n2095_n4160# m4_n33805_n4160# m4_n20315_n4260# m4_2435_n4160# m4_29515_n4260#
+ m4_n6725_n4260# m4_n38435_n4260# m4_25085_n4160# m4_n20215_n4160# m4_15925_n4260#
X0 m4_n42865_n4160# m4_n42965_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X1 m4_n38335_n4160# m4_n38435_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X2 m4_n33805_n4160# m4_n33905_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X3 m4_n29275_n4160# m4_n29375_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X4 m4_n24745_n4160# m4_n24845_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X5 m4_n20215_n4160# m4_n20315_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X6 m4_n15685_n4160# m4_n15785_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X7 m4_n11155_n4160# m4_n11255_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X8 m4_n6625_n4160# m4_n6725_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X9 m4_n2095_n4160# m4_n2195_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X10 m4_2435_n4160# m4_2335_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X11 m4_6965_n4160# m4_6865_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X12 m4_11495_n4160# m4_11395_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X13 m4_16025_n4160# m4_15925_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X14 m4_20555_n4160# m4_20455_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X15 m4_25085_n4160# m4_24985_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X16 m4_29615_n4160# m4_29515_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X17 m4_34145_n4160# m4_34045_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X18 m4_38675_n4160# m4_38575_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X19 m4_n42865_n4160# m4_n42965_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X20 m4_n38335_n4160# m4_n38435_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X21 m4_n33805_n4160# m4_n33905_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X22 m4_n29275_n4160# m4_n29375_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X23 m4_n24745_n4160# m4_n24845_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X24 m4_n20215_n4160# m4_n20315_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X25 m4_n15685_n4160# m4_n15785_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X26 m4_n11155_n4160# m4_n11255_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X27 m4_n6625_n4160# m4_n6725_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X28 m4_n2095_n4160# m4_n2195_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X29 m4_2435_n4160# m4_2335_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X30 m4_6965_n4160# m4_6865_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X31 m4_11495_n4160# m4_11395_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X32 m4_16025_n4160# m4_15925_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X33 m4_20555_n4160# m4_20455_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X34 m4_25085_n4160# m4_24985_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X35 m4_29615_n4160# m4_29515_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X36 m4_34145_n4160# m4_34045_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X37 m4_38675_n4160# m4_38575_n4260# w_n1073741817_n1073741817# cmm5t p=80u a=400p
.ends

* Black-box entry subcircuit for AMUX4_3V abstract view
.subckt AMUX4_3V AIN1 AIN2 AIN3 AIN4 AOUT SEL[0] SEL[1] VDD1V8 VDD3V3 VSSA
.ends

* Black-box entry subcircuit for XSPRAM_1024X32_M8P abstract view
.subckt XSPRAM_1024X32_M8P A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] CEn CLK
+ D[0] D[10] D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[1] D[20] D[21]
+ D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[2] D[30] D[31] D[3] D[4] D[5]
+ D[6] D[7] D[8] D[9] OEn Q[0] Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18]
+ Q[19] Q[1] Q[20] Q[21] Q[22] Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[2] Q[30]
+ Q[31] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] RDY VDD18M VSSM WEn
.ends

* Black-box entry subcircuit for abgpc01_3v3 abstract view
.subckt abgpc01_3v3 VDDA VSSA EN VBGVTN VBGP
.ends

* Black-box entry subcircuit for acmpc01_3v3 abstract view
.subckt acmpc01_3v3 IBN INP INN EN OUT VDDA VSSA
.ends

* Black-box entry subcircuit for acsoc01_3v3 abstract view
.subckt acsoc01_3v3 VDDA VSSA EN CS2_200N CS1_200N CS0_200N CS3_200N
.ends

* Black-box entry subcircuit for arcoc01_3v3 abstract view
.subckt arcoc01_3v3 EN CLK VDDA VSSA
.ends

* Black-box entry subcircuit for aporc02_3v3 abstract view
.subckt aporc02_3v3 POR PORB VDDA VSSA
.ends

.subckt cmm5t_qurpk0 m4_70_n10580# m4_18290_n10480# m4_n4360_n10480# m4_13660_n10580#
+ m4_n22480_n10480# m4_n18050_n10580# m4_4700_n10480# w_n1073741817_n1073741817# m4_13760_n10480#
+ m4_n17950_n10480# m4_n8990_n10580# m4_n13520_n10580# m4_9130_n10580# m4_n8890_n10480#
+ m4_170_n10480# m4_18190_n10580# m4_n13420_n10480# m4_n4460_n10580# m4_n22580_n10580#
+ m4_9230_n10480# m4_4600_n10580#
X0 m4_n22480_n10480# m4_n22580_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X1 m4_n17950_n10480# m4_n18050_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X2 m4_n13420_n10480# m4_n13520_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X3 m4_n8890_n10480# m4_n8990_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X4 m4_n4360_n10480# m4_n4460_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X5 m4_170_n10480# m4_70_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X6 m4_4700_n10480# m4_4600_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X7 m4_9230_n10480# m4_9130_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X8 m4_13760_n10480# m4_13660_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X9 m4_18290_n10480# m4_18190_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X10 m4_n22480_n10480# m4_n22580_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X11 m4_n17950_n10480# m4_n18050_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X12 m4_n13420_n10480# m4_n13520_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X13 m4_n8890_n10480# m4_n8990_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X14 m4_n4360_n10480# m4_n4460_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X15 m4_170_n10480# m4_70_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X16 m4_4700_n10480# m4_4600_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X17 m4_9230_n10480# m4_9130_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X18 m4_13760_n10480# m4_13660_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X19 m4_18290_n10480# m4_18190_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X20 m4_n22480_n10480# m4_n22580_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X21 m4_n17950_n10480# m4_n18050_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X22 m4_n13420_n10480# m4_n13520_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X23 m4_n8890_n10480# m4_n8990_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X24 m4_n4360_n10480# m4_n4460_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X25 m4_170_n10480# m4_70_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X26 m4_4700_n10480# m4_4600_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X27 m4_9230_n10480# m4_9130_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X28 m4_13760_n10480# m4_13660_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X29 m4_18290_n10480# m4_18190_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X30 m4_n22480_n10480# m4_n22580_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X31 m4_n17950_n10480# m4_n18050_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X32 m4_n13420_n10480# m4_n13520_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X33 m4_n8890_n10480# m4_n8990_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X34 m4_n4360_n10480# m4_n4460_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X35 m4_170_n10480# m4_70_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X36 m4_4700_n10480# m4_4600_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X37 m4_9230_n10480# m4_9130_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X38 m4_13760_n10480# m4_13660_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X39 m4_18290_n10480# m4_18190_n10580# w_n1073741817_n1073741817# cmm5t p=90u a=500p
.ends

* Black-box entry subcircuit for raven_spi abstract view
.subckt raven_spi vdd3 gnd RST SCK SDI CSB trap mask_rev_in<0> mask_rev_in<1> mask_rev_in<2>
+ mask_rev_in<3> SDO sdo_enb xtal_ena reg_ena pll_vco_ena pll_cp_ena pll_bias_ena
+ pll_trim<0> pll_trim<1> pll_trim<2> pll_trim<3> pll_bypass irq reset mfgr_id<0>
+ mfgr_id<1> mfgr_id<2> mfgr_id<3> mfgr_id<4> mfgr_id<5> mfgr_id<6> mfgr_id<7> mfgr_id<8>
+ mfgr_id<9> mfgr_id<10> mfgr_id<11> prod_id<0> prod_id<1> prod_id<2> prod_id<3> prod_id<4>
+ prod_id<5> prod_id<6> prod_id<7> mask_rev<0> mask_rev<1> mask_rev<2> mask_rev<3>
.ends

* Black-box entry subcircuit for LS_3VX2 abstract view
.subckt LS_3VX2 VDD1V8 VSSA VDD3V3 A Q
.ends

* Black-box entry subcircuit for BU_3VX2 abstract view
.subckt BU_3VX2 A Q gnd vdd3
.ends

.subckt cmm5t_x3bss8 m4_n11155_n6160# m4_34145_n6160# m4_n29275_n6160# m4_n15785_n6260#
+ m4_24985_n6260# m4_n33905_n6260# m4_n2195_n6260# m4_20555_n6160# m4_6865_n6260#
+ m4_n15685_n6160# m4_11395_n6260# w_n1073741817_n1073741817# m4_n33805_n6160# m4_n2095_n6160#
+ m4_2435_n6160# m4_29515_n6260# m4_n20315_n6260# m4_n38435_n6260# m4_n6725_n6260#
+ m4_25085_n6160# m4_n20215_n6160# m4_15925_n6260# m4_n38335_n6160# m4_n6625_n6160#
+ m4_n24845_n6260# m4_6965_n6160# m4_34045_n6260# m4_11495_n6160# m4_29615_n6160#
+ m4_n24745_n6160# m4_20455_n6260# m4_n11255_n6260# m4_n29375_n6260# m4_16025_n6160#
+ m4_2335_n6260#
X0 m4_n38335_n6160# m4_n38435_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X1 m4_n33805_n6160# m4_n33905_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X2 m4_n29275_n6160# m4_n29375_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X3 m4_n24745_n6160# m4_n24845_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X4 m4_n20215_n6160# m4_n20315_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X5 m4_n15685_n6160# m4_n15785_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X6 m4_n11155_n6160# m4_n11255_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X7 m4_n6625_n6160# m4_n6725_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X8 m4_n2095_n6160# m4_n2195_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X9 m4_2435_n6160# m4_2335_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X10 m4_6965_n6160# m4_6865_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X11 m4_11495_n6160# m4_11395_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X12 m4_16025_n6160# m4_15925_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X13 m4_20555_n6160# m4_20455_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X14 m4_25085_n6160# m4_24985_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X15 m4_29615_n6160# m4_29515_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X16 m4_34145_n6160# m4_34045_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X17 m4_n38335_n6160# m4_n38435_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X18 m4_n33805_n6160# m4_n33905_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X19 m4_n29275_n6160# m4_n29375_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X20 m4_n24745_n6160# m4_n24845_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X21 m4_n20215_n6160# m4_n20315_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X22 m4_n15685_n6160# m4_n15785_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X23 m4_n11155_n6160# m4_n11255_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X24 m4_n6625_n6160# m4_n6725_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X25 m4_n2095_n6160# m4_n2195_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X26 m4_2435_n6160# m4_2335_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X27 m4_6965_n6160# m4_6865_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X28 m4_11495_n6160# m4_11395_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X29 m4_16025_n6160# m4_15925_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X30 m4_20555_n6160# m4_20455_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X31 m4_25085_n6160# m4_24985_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X32 m4_29615_n6160# m4_29515_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X33 m4_34145_n6160# m4_34045_n6260# w_n1073741817_n1073741817# cmm5t p=100u a=600p
.ends

* Black-box entry subcircuit for atmpc01_3v3 abstract view
.subckt atmpc01_3v3 OVT EN VSSA VDDA
.ends

* Black-box entry subcircuit for aopac01_3v3 abstract view
.subckt aopac01_3v3 EN INP INN OUT IB VDDA VSSA
.ends

* Black-box entry subcircuit for acsoc02_3v3 abstract view
.subckt acsoc02_3v3 CS_2U CS_4U EN CS_1U CS_8U VSSA VDDA
.ends

.subckt cmm5t_t9d9xe m4_n2595_n17120# w_n1073741817_n1073741817# m4_n2695_n17220#
X0 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X1 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X2 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X3 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X4 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X5 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X6 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X7 m4_n2595_n17120# m4_n2695_n17220# w_n1073741817_n1073741817# cmm5t p=90u a=500p
.ends

* Black-box entry subcircuit for AMUX2_3V abstract view
.subckt AMUX2_3V AIN1 AIN2 AOUT SEL VDD1V8 VDD3V3 VSSA
.ends

* Black-box entry subcircuit for adacc01_3v3 abstract view
.subckt adacc01_3v3 OUT VSSA VDDA D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0>
+ EN VSS VREFH VREFL VDD
.ends

* Black-box entry subcircuit for raven_soc abstract view
.subckt raven_soc vdd gnd pll_clk ext_clk ext_clk_sel ext_reset reset ram_rdata<0>
+ ram_rdata<1> ram_rdata<2> ram_rdata<3> ram_rdata<4> ram_rdata<5> ram_rdata<6> ram_rdata<7>
+ ram_rdata<8> ram_rdata<9> ram_rdata<10> ram_rdata<11> ram_rdata<12> ram_rdata<13>
+ ram_rdata<14> ram_rdata<15> ram_rdata<16> ram_rdata<17> ram_rdata<18> ram_rdata<19>
+ ram_rdata<20> ram_rdata<21> ram_rdata<22> ram_rdata<23> ram_rdata<24> ram_rdata<25>
+ ram_rdata<26> ram_rdata<27> ram_rdata<28> ram_rdata<29> ram_rdata<30> ram_rdata<31>
+ gpio_in<0> gpio_in<1> gpio_in<2> gpio_in<3> gpio_in<4> gpio_in<5> gpio_in<6> gpio_in<7>
+ gpio_in<8> gpio_in<9> gpio_in<10> gpio_in<11> gpio_in<12> gpio_in<13> gpio_in<14>
+ gpio_in<15> adc0_data<0> adc0_data<1> adc0_data<2> adc0_data<3> adc0_data<4> adc0_data<5>
+ adc0_data<6> adc0_data<7> adc0_data<8> adc0_data<9> adc0_done adc1_data<0> adc1_data<1>
+ adc1_data<2> adc1_data<3> adc1_data<4> adc1_data<5> adc1_data<6> adc1_data<7> adc1_data<8>
+ adc1_data<9> adc1_done overtemp rcosc_in xtal_in comp_in spi_sck spi_ro_config<0>
+ spi_ro_config<1> spi_ro_config<2> spi_ro_config<3> spi_ro_config<4> spi_ro_config<5>
+ spi_ro_config<6> spi_ro_config<7> spi_ro_xtal_ena spi_ro_reg_ena spi_ro_pll_cp_ena
+ spi_ro_pll_vco_ena spi_ro_pll_bias_ena spi_ro_pll_trim<0> spi_ro_pll_trim<1> spi_ro_pll_trim<2>
+ spi_ro_pll_trim<3> spi_ro_mfgr_id<0> spi_ro_mfgr_id<1> spi_ro_mfgr_id<2> spi_ro_mfgr_id<3>
+ spi_ro_mfgr_id<4> spi_ro_mfgr_id<5> spi_ro_mfgr_id<6> spi_ro_mfgr_id<7> spi_ro_mfgr_id<8>
+ spi_ro_mfgr_id<9> spi_ro_mfgr_id<10> spi_ro_mfgr_id<11> spi_ro_prod_id<0> spi_ro_prod_id<1>
+ spi_ro_prod_id<2> spi_ro_prod_id<3> spi_ro_prod_id<4> spi_ro_prod_id<5> spi_ro_prod_id<6>
+ spi_ro_prod_id<7> spi_ro_mask_rev<0> spi_ro_mask_rev<1> spi_ro_mask_rev<2> spi_ro_mask_rev<3>
+ ser_rx irq_pin irq_spi flash_io0_di flash_io1_di flash_io2_di flash_io3_di ram_wenb
+ ram_addr<0> ram_addr<1> ram_addr<2> ram_addr<3> ram_addr<4> ram_addr<5> ram_addr<6>
+ ram_addr<7> ram_addr<8> ram_addr<9> ram_wdata<0> ram_wdata<1> ram_wdata<2> ram_wdata<3>
+ ram_wdata<4> ram_wdata<5> ram_wdata<6> ram_wdata<7> ram_wdata<8> ram_wdata<9> ram_wdata<10>
+ ram_wdata<11> ram_wdata<12> ram_wdata<13> ram_wdata<14> ram_wdata<15> ram_wdata<16>
+ ram_wdata<17> ram_wdata<18> ram_wdata<19> ram_wdata<20> ram_wdata<21> ram_wdata<22>
+ ram_wdata<23> ram_wdata<24> ram_wdata<25> ram_wdata<26> ram_wdata<27> ram_wdata<28>
+ ram_wdata<29> ram_wdata<30> ram_wdata<31> gpio_out<0> gpio_out<1> gpio_out<2> gpio_out<3>
+ gpio_out<4> gpio_out<5> gpio_out<6> gpio_out<7> gpio_out<8> gpio_out<9> gpio_out<10>
+ gpio_out<11> gpio_out<12> gpio_out<13> gpio_out<14> gpio_out<15> gpio_pullup<0>
+ gpio_pullup<1> gpio_pullup<2> gpio_pullup<3> gpio_pullup<4> gpio_pullup<5> gpio_pullup<6>
+ gpio_pullup<7> gpio_pullup<8> gpio_pullup<9> gpio_pullup<10> gpio_pullup<11> gpio_pullup<12>
+ gpio_pullup<13> gpio_pullup<14> gpio_pullup<15> gpio_pulldown<0> gpio_pulldown<1>
+ gpio_pulldown<2> gpio_pulldown<3> gpio_pulldown<4> gpio_pulldown<5> gpio_pulldown<6>
+ gpio_pulldown<7> gpio_pulldown<8> gpio_pulldown<9> gpio_pulldown<10> gpio_pulldown<11>
+ gpio_pulldown<12> gpio_pulldown<13> gpio_pulldown<14> gpio_pulldown<15> gpio_outenb<0>
+ gpio_outenb<1> gpio_outenb<2> gpio_outenb<3> gpio_outenb<4> gpio_outenb<5> gpio_outenb<6>
+ gpio_outenb<7> gpio_outenb<8> gpio_outenb<9> gpio_outenb<10> gpio_outenb<11> gpio_outenb<12>
+ gpio_outenb<13> gpio_outenb<14> gpio_outenb<15> adc0_ena adc0_convert adc0_clk adc0_inputsrc<0>
+ adc0_inputsrc<1> adc1_ena adc1_convert adc1_clk adc1_inputsrc<0> adc1_inputsrc<1>
+ dac_ena dac_value<0> dac_value<1> dac_value<2> dac_value<3> dac_value<4> dac_value<5>
+ dac_value<6> dac_value<7> dac_value<8> dac_value<9> analog_out_sel opamp_ena opamp_bias_ena
+ bg_ena comp_ena comp_ninputsrc<0> comp_ninputsrc<1> comp_pinputsrc<0> comp_pinputsrc<1>
+ rcosc_ena overtemp_ena ser_tx trap flash_csb flash_clk flash_io0_oeb flash_io1_oeb
+ flash_io2_oeb flash_io3_oeb flash_io0_do flash_io1_do flash_io2_do flash_io3_do
.ends

.subckt cmm5t_956f8u m4_6865_n3100# m4_n2095_n3000# m4_2435_n3000# m4_n6725_n3100#
+ w_n1073741817_n1073741817# m4_n6625_n3000# m4_6965_n3000# m4_n11255_n3100# m4_2335_n3100#
+ m4_n11155_n3000# m4_n2195_n3100#
X0 m4_n11155_n3000# m4_n11255_n3100# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X1 m4_n6625_n3000# m4_n6725_n3100# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X2 m4_n2095_n3000# m4_n2195_n3100# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X3 m4_2435_n3000# m4_2335_n3100# w_n1073741817_n1073741817# cmm5t p=100u a=600p
X4 m4_6965_n3000# m4_6865_n3100# w_n1073741817_n1073741817# cmm5t p=100u a=600p
.ends

* Black-box entry subcircuit for aadcc01_3v3 abstract view
.subckt aadcc01_3v3 VDD EOC EN START CLK D<0> D<1> D<2> D<3> D<4> D<5> D<6> D<7> D<8>
+ D<9> VIN VREFH VREFL VSSA VDDA VSS
.ends

.subckt cmm5t_wetxca m4_n18050_n7920# m4_n4460_n7920# m4_9130_n7920# m4_n17950_n7820#
+ m4_13660_n7920# m4_n4360_n7820# m4_4700_n7820# w_n1073741817_n1073741817# m4_n8990_n7920#
+ m4_n8890_n7820# m4_170_n7820# m4_9230_n7820# m4_70_n7920# m4_13760_n7820# m4_n13520_n7920#
+ m4_4600_n7920# m4_n13420_n7820#
X0 m4_n17950_n7820# m4_n18050_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X1 m4_n13420_n7820# m4_n13520_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X2 m4_n8890_n7820# m4_n8990_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X3 m4_n4360_n7820# m4_n4460_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X4 m4_170_n7820# m4_70_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X5 m4_4700_n7820# m4_4600_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X6 m4_9230_n7820# m4_9130_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X7 m4_13760_n7820# m4_13660_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X8 m4_n17950_n7820# m4_n18050_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X9 m4_n13420_n7820# m4_n13520_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X10 m4_n8890_n7820# m4_n8990_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X11 m4_n4360_n7820# m4_n4460_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X12 m4_170_n7820# m4_70_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X13 m4_4700_n7820# m4_4600_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X14 m4_9230_n7820# m4_9130_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X15 m4_13760_n7820# m4_13660_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X16 m4_n17950_n7820# m4_n18050_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X17 m4_n13420_n7820# m4_n13520_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X18 m4_n8890_n7820# m4_n8990_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X19 m4_n4360_n7820# m4_n4460_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X20 m4_170_n7820# m4_70_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X21 m4_4700_n7820# m4_4600_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X22 m4_9230_n7820# m4_9130_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
X23 m4_13760_n7820# m4_13660_n7920# w_n1073741817_n1073741817# cmm5t p=90u a=500p
.ends

* Black-box entry subcircuit for IN_3VX2 abstract view
.subckt IN_3VX2 A Q gnd vdd3
.ends

.subckt cmm5t_zs6qdf m4_n4360_n9680# m4_4700_n9680# m4_n8990_n9780# m4_n8890_n9680#
+ m4_170_n9680# w_n1073741817_n1073741817# m4_70_n9780# m4_4600_n9780# m4_n4460_n9780#
X0 m4_n8890_n9680# m4_n8990_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X1 m4_n4360_n9680# m4_n4460_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X2 m4_170_n9680# m4_70_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X3 m4_4700_n9680# m4_4600_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X4 m4_n8890_n9680# m4_n8990_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X5 m4_n4360_n9680# m4_n4460_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X6 m4_170_n9680# m4_70_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X7 m4_4700_n9680# m4_4600_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X8 m4_n8890_n9680# m4_n8990_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X9 m4_n4360_n9680# m4_n4460_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X10 m4_170_n9680# m4_70_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X11 m4_4700_n9680# m4_4600_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X12 m4_n8890_n9680# m4_n8990_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X13 m4_n4360_n9680# m4_n4460_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X14 m4_170_n9680# m4_70_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
X15 m4_4700_n9680# m4_4600_n9780# w_n1073741817_n1073741817# cmm5t p=86u a=460p
.ends

.subckt cmm5t_hhmkxg m4_18290_n2000# m4_4600_n2100# m4_n13420_n2000# m4_n18050_n2100#
+ m4_n4460_n2100# m4_22820_n2000# w_n1073741817_n1073741817# m4_n17950_n2000# m4_9130_n2100#
+ m4_13660_n2100# m4_n4360_n2000# m4_4700_n2000# m4_n22580_n2100# m4_n8990_n2100#
+ m4_n22480_n2000# m4_18190_n2100# m4_n8890_n2000# m4_170_n2000# m4_9230_n2000# m4_n27110_n2100#
+ m4_13760_n2000# m4_70_n2100# m4_n27010_n2000# m4_n13520_n2100# m4_22720_n2100#
X0 m4_n27010_n2000# m4_n27110_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X1 m4_n22480_n2000# m4_n22580_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X2 m4_n17950_n2000# m4_n18050_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X3 m4_n13420_n2000# m4_n13520_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X4 m4_n8890_n2000# m4_n8990_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X5 m4_n4360_n2000# m4_n4460_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X6 m4_170_n2000# m4_70_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X7 m4_4700_n2000# m4_4600_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X8 m4_9230_n2000# m4_9130_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X9 m4_13760_n2000# m4_13660_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X10 m4_18290_n2000# m4_18190_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X11 m4_22820_n2000# m4_22720_n2100# w_n1073741817_n1073741817# cmm5t p=80u a=400p
.ends

* Black-box entry subcircuit for apllc03_1v8 abstract view
.subckt apllc03_1v8 REF B_VCO B_CP VDDD VSSD B<3> B<2> B<1> B<0> VCO_IN CLK VSSA VDDA
+ EN_CP EN_VCO
.ends

.subckt cmm5t_r1lii0 m4_2835_n3100# w_n1073741817_n1073741817# m4_n2695_n3100# m4_n2595_n3000#
+ m4_2935_n3000# m4_n8225_n3100# m4_n8125_n3000#
X0 m4_n8125_n3000# m4_n8225_n3100# w_n1073741817_n1073741817# cmm5t p=110u a=750p
X1 m4_n2595_n3000# m4_n2695_n3100# w_n1073741817_n1073741817# cmm5t p=110u a=750p
X2 m4_2935_n3000# m4_2835_n3100# w_n1073741817_n1073741817# cmm5t p=110u a=750p
.ends

* Black-box entry subcircuit for acsoc04_1v8 abstract view
.subckt acsoc04_1v8 CS1_2u EN VDDA VSSA CS0_1u CS2_4u CS3_8u
.ends

.subckt cmm5t_vk5q8h m4_n8890_n14960# m4_170_n14960# m4_n4460_n15060# m4_4600_n15060#
+ m4_70_n15060# w_n1073741817_n1073741817# m4_n4360_n14960# m4_4700_n14960# m4_n8990_n15060#
X0 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X1 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X2 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X3 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X4 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X5 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X6 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X7 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X8 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X9 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X10 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X11 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X12 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X13 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X14 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X15 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X16 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X17 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X18 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X19 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X20 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X21 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X22 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X23 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X24 m4_n8890_n14960# m4_n8990_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X25 m4_n4360_n14960# m4_n4460_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X26 m4_170_n14960# m4_70_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
X27 m4_4700_n14960# m4_4600_n15060# w_n1073741817_n1073741817# cmm5t p=80u a=400p
.ends

.subckt raven VDD3V3 vdd VSS XCLK SDI SDO CSB SCK ser_tx ser_rx irq gpio[15] gpio[14]
+ gpio[13] gpio[12] gpio[11] gpio[10] gpio[9] gpio[8] gpio[7] gpio[6] gpio[5] gpio[4]
+ gpio[3] gpio[2] gpio[1] gpio[0] flash_csb flash_clk flash_io0 flash_io1 flash_io2
+ flash_io3 adc_high adc_low adc0_in adc1_in analog_out comp_inp comp_inn XI XO adc0_data<5>
Xraven_padframe_0 LOGIC0_3V_4/Q raven_soc_0/gpio_outenb<4> gpio[10] VDD3V3 XCLK comp_inn
+ raven_soc_0/gpio_pulldown<8> VSS raven_soc_0/gpio_in<5> raven_soc_0/gpio_pullup<9>
+ raven_soc_0/gpio_out<2> LOGIC0_3V_4/Q comp_inp SCK gpio[9] raven_soc_0/flash_io2_do
+ LOGIC0_3V_4/Q raven_soc_0/gpio_outenb<1> flash_io0 comp_inp LOGIC0_3V_4/Q LOGIC0_3V_4/Q
+ raven_soc_0/gpio_pulldown<1> raven_soc_0/irq_pin gpio[14] raven_soc_0/gpio_in<13>
+ raven_soc_0/gpio_pullup<0> raven_soc_0/flash_csb raven_soc_0/gpio_pulldown<13> raven_soc_0/gpio_out<10>
+ vdd gpio[2] raven_soc_0/gpio_pullup<14> raven_soc_0/gpio_in<9> VDD3V3 LOGIC0_3V_4/Q
+ raven_soc_0/gpio_out<6> irq LOGIC0_3V_4/Q raven_soc_0/gpio_pulldown<7> raven_soc_0/gpio_pullup<8>
+ raven_soc_0/gpio_in<1> raven_soc_0/gpio_outenb<14> LOGIC0_3V_4/Q raven_soc_0/flash_io1_oeb
+ raven_soc_0/gpio_outenb<7> raven_soc_0/flash_io1_di LOGIC0_3V_4/Q adc_high raven_soc_0/gpio_out<14>
+ raven_spi_0/SDO gpio[6] raven_spi_0/sdo_enb raven_soc_0/gpio_pulldown<12> raven_soc_0/gpio_pullup<1>
+ gnd raven_soc_0/gpio_pullup<13> BU_3VX2_72/A raven_soc_0/gpio_outenb<10> raven_soc_0/gpio_in<4>
+ raven_soc_0/gpio_outenb<3> gnd gpio[11] raven_soc_0/gpio_out<0> SDI raven_soc_0/flash_io3_do
+ raven_soc_0/gpio_pulldown<6> raven_soc_0/gpio_pullup<7> VDD3V3 LOGIC0_3V_4/Q XCLK
+ raven_soc_0/ser_rx raven_soc_0/gpio_in<12> AMUX4_3V_0/AIN1 raven_soc_0/flash_clk
+ VDD3V3 LOGIC0_3V_4/Q raven_soc_0/gpio_in<8> BU_3VX2_31/A gnd LOGIC0_3V_4/Q LOGIC0_3V_4/Q
+ raven_soc_0/gpio_out<5> flash_io1 raven_soc_0/gpio_pulldown<11> raven_soc_0/gpio_pullup<12>
+ gpio[15] gpio[3] raven_soc_0/flash_io0_di LOGIC0_3V_4/Q IN_3VX2_1/A raven_soc_0/gpio_pulldown<5>
+ raven_soc_0/gpio_pullup<6> BU_3VX2_33/A raven_soc_0/gpio_out<13> raven_soc_0/gpio_outenb<13>
+ LOGIC0_3V_4/Q SDO raven_soc_0/flash_io0_oeb raven_soc_0/gpio_outenb<6> raven_soc_0/gpio_out<9>
+ ser_tx analog_out raven_soc_0/gpio_in<3> IN_3VX2_1/Q gpio[7] raven_soc_0/gpio_out<1>
+ raven_soc_0/gpio_pulldown<10> adc1_in raven_soc_0/flash_io1_do raven_soc_0/gpio_pullup<11>
+ raven_soc_0/gpio_outenb<2> LOGIC0_3V_4/Q LOGIC0_3V_4/Q gpio[12] raven_soc_0/gpio_in<11>
+ gpio[0] raven_soc_0/ser_tx raven_soc_0/gpio_pullup<5> raven_soc_0/gpio_pulldown<4>
+ raven_soc_0/gpio_in<7> flash_csb raven_soc_0/gpio_out<4> LOGIC0_3V_4/Q gnd LOGIC0_3V_4/Q
+ AMUX4_3V_1/AIN1 LOGIC0_3V_4/Q VDD3V3 LOGIC0_3V_4/Q raven_soc_0/flash_io2_oeb raven_soc_0/gpio_outenb<9>
+ raven_soc_0/gpio_pullup<10> flash_io3 raven_soc_0/gpio_in<15> VDD3V3 vdd raven_soc_0/gpio_out<12>
+ raven_spi_0/CSB gpio[4] LOGIC0_3V_4/Q IN_3VX2_1/A raven_soc_0/gpio_out<8> flash_clk
+ raven_soc_0/gpio_pulldown<3> raven_soc_0/gpio_pullup<4> raven_soc_0/gpio_outenb<12>
+ raven_soc_0/gpio_in<2> LOGIC0_3V_4/Q raven_soc_0/flash_io2_di flash_io0 vdd raven_soc_0/gpio_outenb<5>
+ raven_soc_0/flash_io0_do flash_io1 AMUX4_3V_4/AIN1 XI adc0_in flash_io2 gpio[8]
+ IN_3VX2_1/Q raven_soc_0/gpio_in<10> flash_io3 raven_soc_0/gpio_in<6> LOGIC0_3V_4/Q
+ raven_soc_0/gpio_outenb<0> LOGIC0_3V_4/Q LOGIC0_3V_4/Q raven_soc_0/gpio_out<3> gpio[13]
+ vdd raven_soc_0/gpio_pullup<3> raven_soc_0/gpio_pulldown<2> gpio[1] raven_soc_0/gpio_pulldown<15>
+ VDD3V3 CSB raven_soc_0/ext_clk raven_soc_0/gpio_in<14> LOGIC0_3V_4/Q raven_spi_0/SDI
+ flash_clk raven_soc_0/gpio_out<11> raven_soc_0/gpio_pulldown<9> raven_soc_0/gpio_outenb<15>
+ gnd LOGIC0_3V_4/Q ser_rx raven_soc_0/gpio_outenb<8> raven_soc_0/flash_io3_oeb LOGIC0_3V_4/Q
+ adc_low raven_soc_0/gpio_out<7> XO flash_io2 gpio[5] raven_soc_0/gpio_in<0> gnd
+ vdd raven_soc_0/flash_io3_di raven_soc_0/gpio_pulldown<0> VDD3V3 raven_soc_0/gpio_pulldown<14>
+ raven_soc_0/gpio_pullup<15> flash_csb raven_soc_0/gpio_pullup<2> VDD3V3 raven_soc_0/gpio_outenb<11>
+ raven_soc_0/gpio_out<15> raven_padframe
XLOGIC0_3V_4 LOGIC0_3V_4/Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_3 LOGIC0_3V_3/Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_2 LOGIC0_3V_2/Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_1 LOGIC0_3V_1/Q gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_0 LOGIC0_3V_0/Q gnd VDD3V3 LOGIC0_3V
XLOGIC1_3V_3 LOGIC1_3V_3/Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_2 LOGIC1_3V_2/Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_1 LOGIC1_3V_1/Q gnd VDD3V3 LOGIC1_3V
XLOGIC1_3V_0 LOGIC1_3V_0/Q gnd VDD3V3 LOGIC1_3V
Xcmm5t_o8rj96_0 vdd vdd vdd gnd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd gnd vdd gnd
+ vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd gnd vdd gnd gnd gnd vdd
+ vdd gnd cmm5t_o8rj96
XAMUX4_3V_3 comp_inp AMUX4_3V_4/AIN2 AMUX4_3V_4/AIN3 vdd AMUX4_3V_3/AOUT AMUX4_3V_3/SEL[0]
+ AMUX4_3V_3/SEL[1] vdd VDD3V3 gnd AMUX4_3V
XAMUX4_3V_4 AMUX4_3V_4/AIN1 AMUX4_3V_4/AIN2 AMUX4_3V_4/AIN3 vdd AMUX4_3V_4/AOUT AMUX4_3V_4/SEL[0]
+ AMUX4_3V_4/SEL[1] vdd VDD3V3 gnd AMUX4_3V
XXSPRAM_1024X32_M8P_0 raven_soc_0/ram_addr<0> raven_soc_0/ram_addr<1> raven_soc_0/ram_addr<2>
+ raven_soc_0/ram_addr<3> raven_soc_0/ram_addr<4> raven_soc_0/ram_addr<5> raven_soc_0/ram_addr<6>
+ raven_soc_0/ram_addr<7> raven_soc_0/ram_addr<8> raven_soc_0/ram_addr<9> BU_3VX2_0/Q
+ apllc03_1v8_0/CLK raven_soc_0/ram_wdata<0> raven_soc_0/ram_wdata<10> raven_soc_0/ram_wdata<11>
+ raven_soc_0/ram_wdata<12> raven_soc_0/ram_wdata<13> raven_soc_0/ram_wdata<14> raven_soc_0/ram_wdata<15>
+ raven_soc_0/ram_wdata<16> raven_soc_0/ram_wdata<17> raven_soc_0/ram_wdata<18> raven_soc_0/ram_wdata<19>
+ raven_soc_0/ram_wdata<1> raven_soc_0/ram_wdata<20> raven_soc_0/ram_wdata<21> raven_soc_0/ram_wdata<22>
+ raven_soc_0/ram_wdata<23> raven_soc_0/ram_wdata<24> raven_soc_0/ram_wdata<25> raven_soc_0/ram_wdata<26>
+ raven_soc_0/ram_wdata<27> raven_soc_0/ram_wdata<28> raven_soc_0/ram_wdata<29> raven_soc_0/ram_wdata<2>
+ raven_soc_0/ram_wdata<30> raven_soc_0/ram_wdata<31> raven_soc_0/ram_wdata<3> raven_soc_0/ram_wdata<4>
+ raven_soc_0/ram_wdata<5> raven_soc_0/ram_wdata<6> raven_soc_0/ram_wdata<7> raven_soc_0/ram_wdata<8>
+ raven_soc_0/ram_wdata<9> BU_3VX2_0/Q raven_soc_0/ram_rdata<0> raven_soc_0/ram_rdata<10>
+ raven_soc_0/ram_rdata<11> raven_soc_0/ram_rdata<12> raven_soc_0/ram_rdata<13> raven_soc_0/ram_rdata<14>
+ raven_soc_0/ram_rdata<15> raven_soc_0/ram_rdata<16> raven_soc_0/ram_rdata<17> raven_soc_0/ram_rdata<18>
+ raven_soc_0/ram_rdata<19> raven_soc_0/ram_rdata<1> raven_soc_0/ram_rdata<20> raven_soc_0/ram_rdata<21>
+ raven_soc_0/ram_rdata<22> raven_soc_0/ram_rdata<23> raven_soc_0/ram_rdata<24> raven_soc_0/ram_rdata<25>
+ raven_soc_0/ram_rdata<26> raven_soc_0/ram_rdata<27> raven_soc_0/ram_rdata<28> raven_soc_0/ram_rdata<29>
+ raven_soc_0/ram_rdata<2> raven_soc_0/ram_rdata<30> raven_soc_0/ram_rdata<31> raven_soc_0/ram_rdata<3>
+ raven_soc_0/ram_rdata<4> raven_soc_0/ram_rdata<5> raven_soc_0/ram_rdata<6> raven_soc_0/ram_rdata<7>
+ raven_soc_0/ram_rdata<8> raven_soc_0/ram_rdata<9> XSPRAM_1024X32_M8P_0/RDY vdd gnd
+ raven_soc_0/ram_wenb XSPRAM_1024X32_M8P
Xabgpc01_3v3_0 VDD3V3 gnd LS_3VX2_18/Q abgpc01_3v3_0/VBGVTN AMUX4_3V_4/AIN3 abgpc01_3v3
Xacmpc01_3v3_0 acmpc01_3v3_0/IBN AMUX4_3V_3/AOUT AMUX4_3V_4/AOUT LS_3VX2_23/Q BU_3VX2_32/A
+ VDD3V3 gnd acmpc01_3v3
Xacsoc01_3v3_0 VDD3V3 gnd LS_3VX2_23/Q acsoc01_3v3_0/CS2_200N acmpc01_3v3_0/IBN acmpc01_3v3_0/IBN
+ acsoc01_3v3_0/CS3_200N acsoc01_3v3
Xarcoc01_3v3_0 LS_3VX2_2/Q BU_3VX2_1/A VDD3V3 gnd arcoc01_3v3
Xaporc02_3v3_0 BU_3VX2_0/A aporc02_3v3_0/PORB VDD3V3 gnd aporc02_3v3
Xcmm5t_qurpk0_0 vdd VDD3V3 VDD3V3 vdd VDD3V3 vdd VDD3V3 gnd VDD3V3 VDD3V3 vdd vdd
+ vdd VDD3V3 VDD3V3 vdd VDD3V3 vdd vdd VDD3V3 vdd cmm5t_qurpk0
Xraven_spi_0 VDD3V3 gnd BU_3VX2_0/A BU_3VX2_33/A raven_spi_0/SDI raven_spi_0/CSB LS_3VX2_3/Q
+ LOGIC0_3V_0/Q LOGIC0_3V_1/Q LOGIC0_3V_2/Q LOGIC0_3V_3/Q raven_spi_0/SDO raven_spi_0/sdo_enb
+ BU_3VX2_31/A IN_3VX2_1/A BU_3VX2_28/A BU_3VX2_29/A BU_3VX2_27/A BU_3VX2_26/A BU_3VX2_25/A
+ BU_3VX2_24/A BU_3VX2_23/A BU_3VX2_40/A BU_3VX2_71/A BU_3VX2_63/A BU_3VX2_22/A BU_3VX2_21/A
+ BU_3VX2_20/A BU_3VX2_19/A BU_3VX2_18/A BU_3VX2_17/A BU_3VX2_16/A BU_3VX2_15/A BU_3VX2_14/A
+ BU_3VX2_13/A BU_3VX2_12/A BU_3VX2_11/A BU_3VX2_10/A BU_3VX2_9/A BU_3VX2_8/A BU_3VX2_7/A
+ BU_3VX2_6/A BU_3VX2_5/A BU_3VX2_4/A BU_3VX2_3/A BU_3VX2_2/A BU_3VX2_37/A BU_3VX2_38/A
+ BU_3VX2_35/A raven_spi
XLS_3VX2_18 vdd gnd VDD3V3 LS_3VX2_18/A LS_3VX2_18/Q LS_3VX2
XLS_3VX2_23 vdd gnd VDD3V3 LS_3VX2_23/A LS_3VX2_23/Q LS_3VX2
XLS_3VX2_2 vdd gnd VDD3V3 LS_3VX2_2/A LS_3VX2_2/Q LS_3VX2
XBU_3VX2_70 BU_3VX2_70/A BU_3VX2_70/Q gnd vdd BU_3VX2
XBU_3VX2_69 BU_3VX2_69/A BU_3VX2_69/Q gnd vdd BU_3VX2
XBU_3VX2_68 BU_3VX2_68/A BU_3VX2_68/Q gnd vdd BU_3VX2
XBU_3VX2_67 BU_3VX2_67/A BU_3VX2_67/Q gnd vdd BU_3VX2
XBU_3VX2_66 BU_3VX2_66/A BU_3VX2_66/Q gnd vdd BU_3VX2
XBU_3VX2_65 BU_3VX2_65/A BU_3VX2_65/Q gnd vdd BU_3VX2
XBU_3VX2_64 BU_3VX2_64/A BU_3VX2_64/Q gnd vdd BU_3VX2
XBU_3VX2_36 BU_3VX2_36/A BU_3VX2_36/Q gnd vdd BU_3VX2
XBU_3VX2_1 BU_3VX2_1/A BU_3VX2_1/Q gnd vdd BU_3VX2
XBU_3VX2_33 BU_3VX2_33/A BU_3VX2_33/Q gnd vdd BU_3VX2
XBU_3VX2_32 BU_3VX2_32/A BU_3VX2_32/Q gnd vdd BU_3VX2
XLOGIC0_3V_12 BU_3VX2_70/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_11 BU_3VX2_69/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_10 BU_3VX2_68/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_9 BU_3VX2_67/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_8 BU_3VX2_66/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_7 BU_3VX2_65/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_6 BU_3VX2_64/A gnd VDD3V3 LOGIC0_3V
XLOGIC0_3V_5 BU_3VX2_36/A gnd VDD3V3 LOGIC0_3V
XBU_3VX2_0 BU_3VX2_0/A BU_3VX2_0/Q gnd vdd BU_3VX2
XBU_3VX2_31 BU_3VX2_31/A BU_3VX2_31/Q gnd vdd BU_3VX2
XBU_3VX2_30 IN_3VX2_1/A BU_3VX2_30/Q gnd vdd BU_3VX2
XBU_3VX2_29 BU_3VX2_29/A BU_3VX2_29/Q gnd vdd BU_3VX2
XBU_3VX2_28 BU_3VX2_28/A BU_3VX2_28/Q gnd vdd BU_3VX2
XBU_3VX2_27 BU_3VX2_27/A BU_3VX2_27/Q gnd vdd BU_3VX2
XBU_3VX2_26 BU_3VX2_26/A BU_3VX2_26/Q gnd vdd BU_3VX2
XBU_3VX2_25 BU_3VX2_25/A BU_3VX2_25/Q gnd vdd BU_3VX2
XBU_3VX2_24 BU_3VX2_24/A BU_3VX2_24/Q gnd vdd BU_3VX2
XBU_3VX2_23 BU_3VX2_23/A BU_3VX2_23/Q gnd vdd BU_3VX2
XBU_3VX2_22 BU_3VX2_22/A BU_3VX2_22/Q gnd vdd BU_3VX2
XBU_3VX2_21 BU_3VX2_21/A BU_3VX2_21/Q gnd vdd BU_3VX2
XBU_3VX2_20 BU_3VX2_20/A BU_3VX2_20/Q gnd vdd BU_3VX2
XBU_3VX2_19 BU_3VX2_19/A BU_3VX2_19/Q gnd vdd BU_3VX2
XBU_3VX2_18 BU_3VX2_18/A BU_3VX2_18/Q gnd vdd BU_3VX2
XBU_3VX2_17 BU_3VX2_17/A BU_3VX2_17/Q gnd vdd BU_3VX2
XBU_3VX2_16 BU_3VX2_16/A BU_3VX2_16/Q gnd vdd BU_3VX2
XBU_3VX2_15 BU_3VX2_15/A BU_3VX2_15/Q gnd vdd BU_3VX2
XBU_3VX2_14 BU_3VX2_14/A BU_3VX2_14/Q gnd vdd BU_3VX2
XBU_3VX2_13 BU_3VX2_13/A BU_3VX2_13/Q gnd vdd BU_3VX2
XBU_3VX2_12 BU_3VX2_12/A BU_3VX2_12/Q gnd vdd BU_3VX2
XBU_3VX2_11 BU_3VX2_11/A BU_3VX2_11/Q gnd vdd BU_3VX2
XBU_3VX2_10 BU_3VX2_10/A BU_3VX2_10/Q gnd vdd BU_3VX2
XBU_3VX2_9 BU_3VX2_9/A BU_3VX2_9/Q gnd vdd BU_3VX2
XBU_3VX2_8 BU_3VX2_8/A BU_3VX2_8/Q gnd vdd BU_3VX2
XBU_3VX2_7 BU_3VX2_7/A BU_3VX2_7/Q gnd vdd BU_3VX2
XBU_3VX2_6 BU_3VX2_6/A BU_3VX2_6/Q gnd vdd BU_3VX2
XBU_3VX2_5 BU_3VX2_5/A BU_3VX2_5/Q gnd vdd BU_3VX2
XBU_3VX2_4 BU_3VX2_4/A BU_3VX2_4/Q gnd vdd BU_3VX2
XBU_3VX2_3 BU_3VX2_3/A BU_3VX2_3/Q gnd vdd BU_3VX2
XBU_3VX2_2 BU_3VX2_2/A BU_3VX2_2/Q gnd vdd BU_3VX2
XBU_3VX2_37 BU_3VX2_37/A BU_3VX2_37/Q gnd vdd BU_3VX2
XBU_3VX2_38 BU_3VX2_38/A BU_3VX2_38/Q gnd vdd BU_3VX2
XBU_3VX2_35 BU_3VX2_35/A BU_3VX2_35/Q gnd vdd BU_3VX2
XBU_3VX2_40 BU_3VX2_40/A BU_3VX2_40/Q gnd vdd BU_3VX2
XBU_3VX2_63 BU_3VX2_63/A BU_3VX2_63/Q gnd vdd BU_3VX2
XBU_3VX2_71 BU_3VX2_71/A BU_3VX2_71/Q gnd vdd BU_3VX2
XLS_3VX2_3 vdd gnd VDD3V3 LS_3VX2_3/A LS_3VX2_3/Q LS_3VX2
Xcmm5t_x3bss8_0 VDD3V3 VDD3V3 VDD3V3 gnd gnd gnd gnd VDD3V3 gnd VDD3V3 gnd gnd VDD3V3
+ VDD3V3 VDD3V3 gnd gnd gnd gnd VDD3V3 VDD3V3 gnd VDD3V3 VDD3V3 gnd VDD3V3 gnd VDD3V3
+ VDD3V3 VDD3V3 gnd gnd gnd VDD3V3 gnd cmm5t_x3bss8
Xatmpc01_3v3_0 BU_3VX2_73/A LS_3VX2_24/Q gnd VDD3V3 atmpc01_3v3
Xaopac01_3v3_0 LS_3VX2_22/Q AMUX2_3V_0/AOUT analog_out analog_out aopac01_3v3_0/IB
+ VDD3V3 gnd aopac01_3v3
Xacsoc02_3v3_0 aopac01_3v3_0/IB acsoc02_3v3_0/CS_4U LS_3VX2_19/Q aopac01_3v3_0/IB
+ acsoc02_3v3_0/CS_8U gnd VDD3V3 acsoc02_3v3
Xcmm5t_t9d9xe_0 gnd gnd vdd cmm5t_t9d9xe
XLS_3VX2_22 vdd gnd VDD3V3 LS_3VX2_22/A LS_3VX2_22/Q LS_3VX2
XLS_3VX2_19 vdd gnd VDD3V3 LS_3VX2_19/A LS_3VX2_19/Q LS_3VX2
XBU_3VX2_73 BU_3VX2_73/A BU_3VX2_73/Q gnd vdd BU_3VX2
XAMUX2_3V_0 AMUX4_3V_4/AIN2 AMUX4_3V_4/AIN3 AMUX2_3V_0/AOUT AMUX2_3V_0/SEL vdd VDD3V3
+ gnd AMUX2_3V
Xadacc01_3v3_0 AMUX4_3V_4/AIN2 gnd VDD3V3 LS_3VX2_13/Q LS_3VX2_8/Q LS_3VX2_12/Q LS_3VX2_7/Q
+ LS_3VX2_11/Q LS_3VX2_6/Q LS_3VX2_10/Q LS_3VX2_5/Q LS_3VX2_9/Q LS_3VX2_4/Q LS_3VX2_14/Q
+ gnd adc_high adc_low VDD3V3 adacc01_3v3
XLS_3VX2_24 vdd gnd VDD3V3 LS_3VX2_24/A LS_3VX2_24/Q LS_3VX2
XLS_3VX2_4 vdd gnd VDD3V3 LS_3VX2_4/A LS_3VX2_4/Q LS_3VX2
XLS_3VX2_5 vdd gnd VDD3V3 LS_3VX2_5/A LS_3VX2_5/Q LS_3VX2
XLS_3VX2_6 vdd gnd VDD3V3 LS_3VX2_6/A LS_3VX2_6/Q LS_3VX2
XLS_3VX2_7 vdd gnd VDD3V3 LS_3VX2_7/A LS_3VX2_7/Q LS_3VX2
XLS_3VX2_8 vdd gnd VDD3V3 LS_3VX2_8/A LS_3VX2_8/Q LS_3VX2
XLS_3VX2_14 vdd gnd VDD3V3 LS_3VX2_14/A LS_3VX2_14/Q LS_3VX2
XLS_3VX2_9 vdd gnd VDD3V3 LS_3VX2_9/A LS_3VX2_9/Q LS_3VX2
XLS_3VX2_10 vdd gnd VDD3V3 LS_3VX2_10/A LS_3VX2_10/Q LS_3VX2
XLS_3VX2_11 vdd gnd VDD3V3 LS_3VX2_11/A LS_3VX2_11/Q LS_3VX2
XLS_3VX2_12 vdd gnd VDD3V3 LS_3VX2_12/A LS_3VX2_12/Q LS_3VX2
XLS_3VX2_13 vdd gnd VDD3V3 LS_3VX2_13/A LS_3VX2_13/Q LS_3VX2
Xraven_soc_0 vdd gnd apllc03_1v8_0/CLK raven_soc_0/ext_clk BU_3VX2_40/Q BU_3VX2_63/Q
+ BU_3VX2_0/Q raven_soc_0/ram_rdata<0> raven_soc_0/ram_rdata<1> raven_soc_0/ram_rdata<2>
+ raven_soc_0/ram_rdata<3> raven_soc_0/ram_rdata<4> raven_soc_0/ram_rdata<5> raven_soc_0/ram_rdata<6>
+ raven_soc_0/ram_rdata<7> raven_soc_0/ram_rdata<8> raven_soc_0/ram_rdata<9> raven_soc_0/ram_rdata<10>
+ raven_soc_0/ram_rdata<11> raven_soc_0/ram_rdata<12> raven_soc_0/ram_rdata<13> raven_soc_0/ram_rdata<14>
+ raven_soc_0/ram_rdata<15> raven_soc_0/ram_rdata<16> raven_soc_0/ram_rdata<17> raven_soc_0/ram_rdata<18>
+ raven_soc_0/ram_rdata<19> raven_soc_0/ram_rdata<20> raven_soc_0/ram_rdata<21> raven_soc_0/ram_rdata<22>
+ raven_soc_0/ram_rdata<23> raven_soc_0/ram_rdata<24> raven_soc_0/ram_rdata<25> raven_soc_0/ram_rdata<26>
+ raven_soc_0/ram_rdata<27> raven_soc_0/ram_rdata<28> raven_soc_0/ram_rdata<29> raven_soc_0/ram_rdata<30>
+ raven_soc_0/ram_rdata<31> raven_soc_0/gpio_in<0> raven_soc_0/gpio_in<1> raven_soc_0/gpio_in<2>
+ raven_soc_0/gpio_in<3> raven_soc_0/gpio_in<4> raven_soc_0/gpio_in<5> raven_soc_0/gpio_in<6>
+ raven_soc_0/gpio_in<7> raven_soc_0/gpio_in<8> raven_soc_0/gpio_in<9> raven_soc_0/gpio_in<10>
+ raven_soc_0/gpio_in<11> raven_soc_0/gpio_in<12> raven_soc_0/gpio_in<13> raven_soc_0/gpio_in<14>
+ raven_soc_0/gpio_in<15> BU_3VX2_43/Q BU_3VX2_44/Q BU_3VX2_45/Q BU_3VX2_46/Q adc0_data<5>
+ BU_3VX2_47/Q BU_3VX2_48/Q BU_3VX2_49/Q BU_3VX2_50/Q BU_3VX2_51/Q BU_3VX2_42/Q BU_3VX2_61/Q
+ BU_3VX2_60/Q BU_3VX2_59/Q BU_3VX2_58/Q BU_3VX2_57/Q BU_3VX2_56/Q BU_3VX2_55/Q BU_3VX2_54/Q
+ BU_3VX2_53/Q BU_3VX2_52/Q BU_3VX2_62/Q BU_3VX2_73/Q BU_3VX2_1/Q BU_3VX2_72/Q BU_3VX2_32/Q
+ BU_3VX2_33/Q BU_3VX2_36/Q BU_3VX2_64/Q BU_3VX2_65/Q BU_3VX2_66/Q BU_3VX2_67/Q BU_3VX2_68/Q
+ BU_3VX2_69/Q BU_3VX2_70/Q BU_3VX2_31/Q BU_3VX2_30/Q BU_3VX2_29/Q BU_3VX2_28/Q BU_3VX2_27/Q
+ BU_3VX2_26/Q BU_3VX2_25/Q BU_3VX2_24/Q BU_3VX2_23/Q BU_3VX2_22/Q BU_3VX2_21/Q BU_3VX2_20/Q
+ BU_3VX2_19/Q BU_3VX2_18/Q BU_3VX2_17/Q BU_3VX2_16/Q BU_3VX2_15/Q BU_3VX2_14/Q BU_3VX2_13/Q
+ BU_3VX2_12/Q BU_3VX2_11/Q BU_3VX2_10/Q BU_3VX2_9/Q BU_3VX2_8/Q BU_3VX2_7/Q BU_3VX2_6/Q
+ BU_3VX2_5/Q BU_3VX2_4/Q BU_3VX2_3/Q BU_3VX2_2/Q BU_3VX2_37/Q BU_3VX2_38/Q BU_3VX2_35/Q
+ raven_soc_0/ser_rx raven_soc_0/irq_pin BU_3VX2_71/Q raven_soc_0/flash_io0_di raven_soc_0/flash_io1_di
+ raven_soc_0/flash_io2_di raven_soc_0/flash_io3_di raven_soc_0/ram_wenb raven_soc_0/ram_addr<0>
+ raven_soc_0/ram_addr<1> raven_soc_0/ram_addr<2> raven_soc_0/ram_addr<3> raven_soc_0/ram_addr<4>
+ raven_soc_0/ram_addr<5> raven_soc_0/ram_addr<6> raven_soc_0/ram_addr<7> raven_soc_0/ram_addr<8>
+ raven_soc_0/ram_addr<9> raven_soc_0/ram_wdata<0> raven_soc_0/ram_wdata<1> raven_soc_0/ram_wdata<2>
+ raven_soc_0/ram_wdata<3> raven_soc_0/ram_wdata<4> raven_soc_0/ram_wdata<5> raven_soc_0/ram_wdata<6>
+ raven_soc_0/ram_wdata<7> raven_soc_0/ram_wdata<8> raven_soc_0/ram_wdata<9> raven_soc_0/ram_wdata<10>
+ raven_soc_0/ram_wdata<11> raven_soc_0/ram_wdata<12> raven_soc_0/ram_wdata<13> raven_soc_0/ram_wdata<14>
+ raven_soc_0/ram_wdata<15> raven_soc_0/ram_wdata<16> raven_soc_0/ram_wdata<17> raven_soc_0/ram_wdata<18>
+ raven_soc_0/ram_wdata<19> raven_soc_0/ram_wdata<20> raven_soc_0/ram_wdata<21> raven_soc_0/ram_wdata<22>
+ raven_soc_0/ram_wdata<23> raven_soc_0/ram_wdata<24> raven_soc_0/ram_wdata<25> raven_soc_0/ram_wdata<26>
+ raven_soc_0/ram_wdata<27> raven_soc_0/ram_wdata<28> raven_soc_0/ram_wdata<29> raven_soc_0/ram_wdata<30>
+ raven_soc_0/ram_wdata<31> raven_soc_0/gpio_out<0> raven_soc_0/gpio_out<1> raven_soc_0/gpio_out<2>
+ raven_soc_0/gpio_out<3> raven_soc_0/gpio_out<4> raven_soc_0/gpio_out<5> raven_soc_0/gpio_out<6>
+ raven_soc_0/gpio_out<7> raven_soc_0/gpio_out<8> raven_soc_0/gpio_out<9> raven_soc_0/gpio_out<10>
+ raven_soc_0/gpio_out<11> raven_soc_0/gpio_out<12> raven_soc_0/gpio_out<13> raven_soc_0/gpio_out<14>
+ raven_soc_0/gpio_out<15> raven_soc_0/gpio_pullup<0> raven_soc_0/gpio_pullup<1> raven_soc_0/gpio_pullup<2>
+ raven_soc_0/gpio_pullup<3> raven_soc_0/gpio_pullup<4> raven_soc_0/gpio_pullup<5>
+ raven_soc_0/gpio_pullup<6> raven_soc_0/gpio_pullup<7> raven_soc_0/gpio_pullup<8>
+ raven_soc_0/gpio_pullup<9> raven_soc_0/gpio_pullup<10> raven_soc_0/gpio_pullup<11>
+ raven_soc_0/gpio_pullup<12> raven_soc_0/gpio_pullup<13> raven_soc_0/gpio_pullup<14>
+ raven_soc_0/gpio_pullup<15> raven_soc_0/gpio_pulldown<0> raven_soc_0/gpio_pulldown<1>
+ raven_soc_0/gpio_pulldown<2> raven_soc_0/gpio_pulldown<3> raven_soc_0/gpio_pulldown<4>
+ raven_soc_0/gpio_pulldown<5> raven_soc_0/gpio_pulldown<6> raven_soc_0/gpio_pulldown<7>
+ raven_soc_0/gpio_pulldown<8> raven_soc_0/gpio_pulldown<9> raven_soc_0/gpio_pulldown<10>
+ raven_soc_0/gpio_pulldown<11> raven_soc_0/gpio_pulldown<12> raven_soc_0/gpio_pulldown<13>
+ raven_soc_0/gpio_pulldown<14> raven_soc_0/gpio_pulldown<15> raven_soc_0/gpio_outenb<0>
+ raven_soc_0/gpio_outenb<1> raven_soc_0/gpio_outenb<2> raven_soc_0/gpio_outenb<3>
+ raven_soc_0/gpio_outenb<4> raven_soc_0/gpio_outenb<5> raven_soc_0/gpio_outenb<6>
+ raven_soc_0/gpio_outenb<7> raven_soc_0/gpio_outenb<8> raven_soc_0/gpio_outenb<9>
+ raven_soc_0/gpio_outenb<10> raven_soc_0/gpio_outenb<11> raven_soc_0/gpio_outenb<12>
+ raven_soc_0/gpio_outenb<13> raven_soc_0/gpio_outenb<14> raven_soc_0/gpio_outenb<15>
+ LS_3VX2_27/A LS_3VX2_21/A LS_3VX2_20/A AMUX4_3V_0/SEL[0] AMUX4_3V_0/SEL[1] LS_3VX2_17/A
+ LS_3VX2_16/A LS_3VX2_15/A AMUX4_3V_1/SEL[0] AMUX4_3V_1/SEL[1] LS_3VX2_14/A LS_3VX2_4/A
+ LS_3VX2_9/A LS_3VX2_5/A LS_3VX2_10/A LS_3VX2_6/A LS_3VX2_11/A LS_3VX2_7/A LS_3VX2_12/A
+ LS_3VX2_8/A LS_3VX2_13/A AMUX2_3V_0/SEL LS_3VX2_22/A LS_3VX2_19/A LS_3VX2_18/A LS_3VX2_23/A
+ AMUX4_3V_4/SEL[0] AMUX4_3V_4/SEL[1] AMUX4_3V_3/SEL[0] AMUX4_3V_3/SEL[1] LS_3VX2_2/A
+ LS_3VX2_24/A raven_soc_0/ser_tx LS_3VX2_3/A raven_soc_0/flash_csb raven_soc_0/flash_clk
+ raven_soc_0/flash_io0_oeb raven_soc_0/flash_io1_oeb raven_soc_0/flash_io2_oeb raven_soc_0/flash_io3_oeb
+ raven_soc_0/flash_io0_do raven_soc_0/flash_io1_do raven_soc_0/flash_io2_do raven_soc_0/flash_io3_do
+ raven_soc
Xcmm5t_956f8u_0 VDD3V3 gnd gnd VDD3V3 gnd gnd gnd VDD3V3 VDD3V3 gnd VDD3V3 cmm5t_956f8u
Xaadcc01_3v3_0 VDD3V3 BU_3VX2_62/A LS_3VX2_17/Q LS_3VX2_16/Q LS_3VX2_15/Q BU_3VX2_61/A
+ BU_3VX2_60/A BU_3VX2_59/A BU_3VX2_58/A BU_3VX2_57/A BU_3VX2_56/A BU_3VX2_55/A BU_3VX2_54/A
+ BU_3VX2_53/A BU_3VX2_52/A AMUX4_3V_1/AOUT adc_high adc_low gnd VDD3V3 gnd aadcc01_3v3
XAMUX4_3V_1 AMUX4_3V_1/AIN1 VDD3V3 AMUX4_3V_4/AIN3 comp_inp AMUX4_3V_1/AOUT AMUX4_3V_1/SEL[0]
+ AMUX4_3V_1/SEL[1] vdd VDD3V3 gnd AMUX4_3V
Xcmm5t_wetxca_0 gnd gnd gnd VDD3V3 gnd VDD3V3 VDD3V3 gnd gnd VDD3V3 VDD3V3 VDD3V3
+ gnd VDD3V3 gnd gnd VDD3V3 cmm5t_wetxca
Xaadcc01_3v3_1 VDD3V3 BU_3VX2_42/A LS_3VX2_27/Q LS_3VX2_21/Q LS_3VX2_20/Q BU_3VX2_43/A
+ BU_3VX2_44/A BU_3VX2_45/A BU_3VX2_46/A BU_3VX2_41/A BU_3VX2_47/A BU_3VX2_48/A BU_3VX2_49/A
+ BU_3VX2_50/A BU_3VX2_51/A AMUX4_3V_0/AOUT adc_high adc_low gnd VDD3V3 gnd aadcc01_3v3
XIN_3VX2_1 IN_3VX2_1/A IN_3VX2_1/Q gnd VDD3V3 IN_3VX2
XAMUX4_3V_0 AMUX4_3V_0/AIN1 vdd AMUX4_3V_4/AIN2 gnd AMUX4_3V_0/AOUT AMUX4_3V_0/SEL[0]
+ AMUX4_3V_0/SEL[1] vdd VDD3V3 gnd AMUX4_3V
XLS_3VX2_17 vdd gnd VDD3V3 LS_3VX2_17/A LS_3VX2_17/Q LS_3VX2
XLS_3VX2_16 vdd gnd VDD3V3 LS_3VX2_16/A LS_3VX2_16/Q LS_3VX2
XLS_3VX2_15 vdd gnd VDD3V3 LS_3VX2_15/A LS_3VX2_15/Q LS_3VX2
XBU_3VX2_62 BU_3VX2_62/A BU_3VX2_62/Q gnd vdd BU_3VX2
XBU_3VX2_61 BU_3VX2_61/A BU_3VX2_61/Q gnd vdd BU_3VX2
XBU_3VX2_60 BU_3VX2_60/A BU_3VX2_60/Q gnd vdd BU_3VX2
XBU_3VX2_59 BU_3VX2_59/A BU_3VX2_59/Q gnd vdd BU_3VX2
XBU_3VX2_58 BU_3VX2_58/A BU_3VX2_58/Q gnd vdd BU_3VX2
XBU_3VX2_57 BU_3VX2_57/A BU_3VX2_57/Q gnd vdd BU_3VX2
XBU_3VX2_56 BU_3VX2_56/A BU_3VX2_56/Q gnd vdd BU_3VX2
XBU_3VX2_55 BU_3VX2_55/A BU_3VX2_55/Q gnd vdd BU_3VX2
XBU_3VX2_54 BU_3VX2_54/A BU_3VX2_54/Q gnd vdd BU_3VX2
XBU_3VX2_53 BU_3VX2_53/A BU_3VX2_53/Q gnd vdd BU_3VX2
XBU_3VX2_52 BU_3VX2_52/A BU_3VX2_52/Q gnd vdd BU_3VX2
Xcmm5t_zs6qdf_0 vdd vdd gnd vdd vdd gnd gnd gnd gnd cmm5t_zs6qdf
Xcmm5t_hhmkxg_0 gnd VDD3V3 gnd VDD3V3 VDD3V3 gnd gnd gnd VDD3V3 VDD3V3 gnd gnd VDD3V3
+ VDD3V3 gnd VDD3V3 gnd gnd gnd VDD3V3 gnd VDD3V3 gnd VDD3V3 VDD3V3 cmm5t_hhmkxg
XLS_3VX2_27 vdd gnd VDD3V3 LS_3VX2_27/A LS_3VX2_27/Q LS_3VX2
XLS_3VX2_21 vdd gnd VDD3V3 LS_3VX2_21/A LS_3VX2_21/Q LS_3VX2
XLS_3VX2_20 vdd gnd VDD3V3 LS_3VX2_20/A LS_3VX2_20/Q LS_3VX2
XBU_3VX2_42 BU_3VX2_42/A BU_3VX2_42/Q gnd vdd BU_3VX2
XBU_3VX2_43 BU_3VX2_43/A BU_3VX2_43/Q gnd vdd BU_3VX2
XBU_3VX2_44 BU_3VX2_44/A BU_3VX2_44/Q gnd vdd BU_3VX2
XBU_3VX2_45 BU_3VX2_45/A BU_3VX2_45/Q gnd vdd BU_3VX2
XBU_3VX2_46 BU_3VX2_46/A BU_3VX2_46/Q gnd vdd BU_3VX2
XBU_3VX2_41 BU_3VX2_41/A adc0_data<5> gnd vdd BU_3VX2
XBU_3VX2_47 BU_3VX2_47/A BU_3VX2_47/Q gnd vdd BU_3VX2
XBU_3VX2_48 BU_3VX2_48/A BU_3VX2_48/Q gnd vdd BU_3VX2
XBU_3VX2_49 BU_3VX2_49/A BU_3VX2_49/Q gnd vdd BU_3VX2
XBU_3VX2_50 BU_3VX2_50/A BU_3VX2_50/Q gnd vdd BU_3VX2
XBU_3VX2_51 BU_3VX2_51/A BU_3VX2_51/Q gnd vdd BU_3VX2
Xapllc03_1v8_0 BU_3VX2_72/Q apllc03_1v8_0/B_VCO apllc03_1v8_0/B_CP vdd gnd BU_3VX2_23/Q
+ BU_3VX2_24/Q BU_3VX2_25/Q BU_3VX2_26/Q apllc03_1v8_0/VCO_IN apllc03_1v8_0/CLK gnd
+ vdd BU_3VX2_29/Q BU_3VX2_28/Q apllc03_1v8
Xcmm5t_r1lii0_0 gnd gnd gnd VDD3V3 VDD3V3 gnd VDD3V3 cmm5t_r1lii0
Xacsoc04_1v8_0 apllc03_1v8_0/B_CP BU_3VX2_27/Q vdd gnd apllc03_1v8_0/B_VCO apllc03_1v8_0/B_VCO
+ apllc03_1v8_0/B_CP acsoc04_1v8
Xcmm5t_vk5q8h_0 VDD3V3 VDD3V3 gnd gnd gnd gnd VDD3V3 VDD3V3 gnd cmm5t_vk5q8h
XBU_3VX2_72 BU_3VX2_72/A BU_3VX2_72/Q gnd vdd BU_3VX2
.ends

